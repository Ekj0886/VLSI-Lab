****  Final Project: Two stage pipeline Two mode 6-bit MAC  ***

*************************************************************
*************************************************************
***************Don't touch settings below********************
*************************************************************
*************************************************************
.lib "umc018.l" L18U18V_TT 
.vec 'MAC6.vec'

.temp 25
.op
.options brief post

***************** parameter ****************************
.global  VDD  GND
.param supply = 1.8v
.param load = 10f
.param tr = 0.2n

***************** voltage source ****************************
Vclk CLK GND pulse(0 supply 0 0.1ns 0.1ns "1*period/2-tr" "period*1")
Vd1 VDD GND supply

***************** top-circuit ****************************
XMAC6   VDD GND CLK ACC[1] ACC[2] ACC[4] ACC[6] ACC[8] ACC[10] ACC[0]
+ ACC[3] ACC[5] ACC[7] ACC[9] ACC[11] MODE OUT[0] OUT[1] OUT[2] OUT[3] OUT[4]
+ OUT[5] OUT[6] OUT[8] OUT[9] OUT[7] OUT[10] OUT[11] OUT[12] A[4] A[5] A[3] A[2]
+ A[0] A[1] B[0] B[1] B[2] B[3] B[4] B[5] MAC6
     
CLOAD01 OUT[0] GND load
CLOAD02 OUT[1] GND load 
CLOAD03 OUT[2] GND load 
CLOAD04 OUT[3] GND load 
CLOAD05 OUT[4] GND load 
CLOAD06 OUT[5] GND load 
CLOAD07 OUT[6] GND load 
CLOAD08 OUT[7] GND load 
CLOAD09 OUT[8] GND load 
CLOAD10 OUT[9] GND load 
CLOAD11 OUT[10] GND load 
CLOAD12 OUT[11] GND load 
CLOAD13 OUT[12] GND load 

***************** Average Power ****************************
.meas tran Iavg avg I(Vd1) from=0ns to='100*period'
.meas Pavg param='abs(Iavg)*supply'

.tran 0.1n '1000*period'

*************************************************************
*************************************************************
***************Don't touch settings above********************
*************************************************************
*************************************************************

***** you can modify clock cycle here, remember synchronize with clock cycle in MAC6.vec ****
.param period = 5n


* File: MAC6_LPE.sp
* Created: Thu Jan 12 23:02:48 2023
* Program "Calibre xRC"
* Version "v2021.1_33.19"
* 
.include "MAC6_LPE.sp.pex"
.subckt MAC6  VDD GND CLK ACC[1] ACC[2] ACC[4] ACC[6] ACC[8] ACC[10] ACC[0]
+ ACC[3] ACC[5] ACC[7] ACC[9] ACC[11] MODE OUT[0] OUT[1] OUT[2] OUT[3] OUT[4]
+ OUT[5] OUT[6] OUT[8] OUT[9] OUT[7] OUT[10] OUT[11] OUT[12] A[4] A[5] A[3] A[2]
+ A[0] A[1] B[0] B[1] B[2] B[3] B[4] B[5]
* 
* B[5]	B[5]
* B[4]	B[4]
* B[3]	B[3]
* B[2]	B[2]
* B[1]	B[1]
* B[0]	B[0]
* A[1]	A[1]
* A[0]	A[0]
* A[2]	A[2]
* A[3]	A[3]
* A[5]	A[5]
* A[4]	A[4]
* OUT[12]	OUT[12]
* OUT[11]	OUT[11]
* OUT[10]	OUT[10]
* OUT[7]	OUT[7]
* OUT[9]	OUT[9]
* OUT[8]	OUT[8]
* OUT[6]	OUT[6]
* OUT[5]	OUT[5]
* OUT[4]	OUT[4]
* OUT[3]	OUT[3]
* OUT[2]	OUT[2]
* OUT[1]	OUT[1]
* OUT[0]	OUT[0]
* MODE	MODE
* ACC[11]	ACC[11]
* ACC[9]	ACC[9]
* ACC[7]	ACC[7]
* ACC[5]	ACC[5]
* ACC[3]	ACC[3]
* ACC[0]	ACC[0]
* ACC[10]	ACC[10]
* ACC[8]	ACC[8]
* ACC[6]	ACC[6]
* ACC[4]	ACC[4]
* ACC[2]	ACC[2]
* ACC[1]	ACC[1]
* CLK	CLK
* GND	GND
* VDD	VDD
mXADDER/Xa000/Xao1/M10 N_XADDER/XA000/XAO1/N004_XADDER/Xa000/Xao1/M10_d
+ N_CIN_XADDER/Xa000/Xao1/M10_g N_GND_XADDER/Xa000/Xao1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXADDER/Xa01/Xrb2/M3 N_XADDER/P0_XADDER/Xa01/Xrb2/M3_d
+ N_XADDER/XA01/XRB2/N002_XADDER/Xa01/Xrb2/M3_g N_GND_XADDER/Xa01/Xrb2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa72/M3 N_OUT1[2]_XADDER/Xa72/M3_d N_XADDER/XA72/N002_XADDER/Xa72/M3_g
+ N_GND_XADDER/Xa72/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa000/Xao1/M9 N_XADDER/XA000/XAO1/N003_XADDER/Xa000/Xao1/M9_d
+ N_XADDER/P0_XADDER/Xa000/Xao1/M9_g
+ N_XADDER/XA000/XAO1/N004_XADDER/Xa000/Xao1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b
+ N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=6.16e-14 PD=1.74e-06 PS=2.8e-07
mXADDER/Xa70/M2 N_XADDER/XA70/N002_XADDER/Xa70/M2_d N_XADDER/P0_XADDER/Xa70/M2_g
+ N_CIN_XADDER/Xa70/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xdffa4/M3 N_XBOOTH/XDFFA4/N0_XBOOTH/Xdffa4/M3_d
+ N_A[4]_XBOOTH/Xdffa4/M3_g N_GND_XBOOTH/Xdffa4/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xdffa5/M3 N_XBOOTH/XDFFA5/N0_XBOOTH/Xdffa5/M3_d
+ N_A[5]_XBOOTH/Xdffa5/M3_g N_GND_XBOOTH/Xdffa5/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xdffa3/M3 N_XBOOTH/XDFFA3/N0_XBOOTH/Xdffa3/M3_d
+ N_A[3]_XBOOTH/Xdffa3/M3_g N_GND_XBOOTH/Xdffa3/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xdffa2/M3 N_XBOOTH/XDFFA2/N0_XBOOTH/Xdffa2/M3_d
+ N_A[2]_XBOOTH/Xdffa2/M3_g N_GND_XBOOTH/Xdffa2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xdffa0/M3 N_XBOOTH/XDFFA0/N0_XBOOTH/Xdffa0/M3_d
+ N_A[0]_XBOOTH/Xdffa0/M3_g N_GND_XBOOTH/Xdffa0/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xdffa1/M3 N_XBOOTH/XDFFA1/N0_XBOOTH/Xdffa1/M3_d
+ N_A[1]_XBOOTH/Xdffa1/M3_g N_GND_XBOOTH/Xdffa1/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa70/M1 N_XADDER/XA70/N002_XADDER/Xa70/M1_d N_CIN_XADDER/Xa70/M1_g
+ N_XADDER/P0_XADDER/Xa70/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=2.332e-13 PD=5.4e-07 PS=1.5e-06
mXADDER/Xa01/Xrb2/M1 N_XADDER/XA01/XRB2/N002_XADDER/Xa01/Xrb2/M1_d
+ N_GND_XADDER/Xa01/Xrb2/M1_g N_S[0]_XADDER/Xa01/Xrb2/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xdffa4/M6 N_XBOOTH/XDFFA4/P002_XBOOTH/Xdffa4/M6_d
+ N_CLK_XBOOTH/Xdffa4/M6_g N_GND_XBOOTH/Xdffa4/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXBOOTH/Xdffa5/M6 N_XBOOTH/XDFFA5/P002_XBOOTH/Xdffa5/M6_d
+ N_CLK_XBOOTH/Xdffa5/M6_g N_GND_XBOOTH/Xdffa5/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXBOOTH/Xdffa3/M6 N_XBOOTH/XDFFA3/P002_XBOOTH/Xdffa3/M6_d
+ N_CLK_XBOOTH/Xdffa3/M6_g N_GND_XBOOTH/Xdffa3/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXBOOTH/Xdffa2/M6 N_XBOOTH/XDFFA2/P002_XBOOTH/Xdffa2/M6_d
+ N_CLK_XBOOTH/Xdffa2/M6_g N_GND_XBOOTH/Xdffa2/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXBOOTH/Xdffa0/M6 N_XBOOTH/XDFFA0/P002_XBOOTH/Xdffa0/M6_d
+ N_CLK_XBOOTH/Xdffa0/M6_g N_GND_XBOOTH/Xdffa0/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXBOOTH/Xdffa1/M6 N_XBOOTH/XDFFA1/P002_XBOOTH/Xdffa1/M6_d
+ N_CLK_XBOOTH/Xdffa1/M6_g N_GND_XBOOTH/Xdffa1/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXADDER/Xa000/Xao1/Xand1/M16 N_XADDER/XA000/OUT1_XADDER/Xa000/Xao1/Xand1/M16_d
+ N_XADDER/XA000/XAO1/N003_XADDER/Xa000/Xao1/Xand1/M16_g
+ N_GND_XADDER/Xa000/Xao1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xdffa4/M5 N_XBOOTH/XDFFA4/N1_XBOOTH/Xdffa4/M5_d
+ N_XBOOTH/XDFFA4/N0_XBOOTH/Xdffa4/M5_g N_XBOOTH/XDFFA4/P002_XBOOTH/Xdffa4/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xdffa5/M5 N_XBOOTH/XDFFA5/N1_XBOOTH/Xdffa5/M5_d
+ N_XBOOTH/XDFFA5/N0_XBOOTH/Xdffa5/M5_g N_XBOOTH/XDFFA5/P002_XBOOTH/Xdffa5/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xdffa3/M5 N_XBOOTH/XDFFA3/N1_XBOOTH/Xdffa3/M5_d
+ N_XBOOTH/XDFFA3/N0_XBOOTH/Xdffa3/M5_g N_XBOOTH/XDFFA3/P002_XBOOTH/Xdffa3/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xdffa2/M5 N_XBOOTH/XDFFA2/N1_XBOOTH/Xdffa2/M5_d
+ N_XBOOTH/XDFFA2/N0_XBOOTH/Xdffa2/M5_g N_XBOOTH/XDFFA2/P002_XBOOTH/Xdffa2/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xdffa0/M5 N_XBOOTH/XDFFA0/N1_XBOOTH/Xdffa0/M5_d
+ N_XBOOTH/XDFFA0/N0_XBOOTH/Xdffa0/M5_g N_XBOOTH/XDFFA0/P002_XBOOTH/Xdffa0/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xdffa1/M5 N_XBOOTH/XDFFA1/N1_XBOOTH/Xdffa1/M5_d
+ N_XBOOTH/XDFFA1/N0_XBOOTH/Xdffa1/M5_g N_XBOOTH/XDFFA1/P002_XBOOTH/Xdffa1/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa01/Xrb2/M2 N_XADDER/XA01/XRB2/N002_XADDER/Xa01/Xrb2/M2_d
+ N_S[0]_XADDER/Xa01/Xrb2/M2_g N_GND_XADDER/Xa01/Xrb2/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXADDER/Xa72/M1 N_XADDER/XA72/N002_XADDER/Xa72/M1_d N_XADDER/P2_XADDER/Xa72/M1_g
+ N_XADDER/GG1_XADDER/Xa72/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=2.332e-13 PD=5.4e-07 PS=1.5e-06
mXACCXOR/X_xor1/M3 N_CACC[1]_XACCXOR/X_xor1/M3_d
+ N_XACCXOR/X_XOR1/N002_XACCXOR/X_xor1/M3_g N_GND_XACCXOR/X_xor1/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor2/M3 N_CACC[2]_XACCXOR/X_xor2/M3_d
+ N_XACCXOR/X_XOR2/N002_XACCXOR/X_xor2/M3_g N_GND_XACCXOR/X_xor2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor4/M3 N_CACC[4]_XACCXOR/X_xor4/M3_d
+ N_XACCXOR/X_XOR4/N002_XACCXOR/X_xor4/M3_g N_GND_XACCXOR/X_xor4/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor6/M3 N_CACC[6]_XACCXOR/X_xor6/M3_d
+ N_XACCXOR/X_XOR6/N002_XACCXOR/X_xor6/M3_g N_GND_XACCXOR/X_xor6/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor8/M3 N_CACC[8]_XACCXOR/X_xor8/M3_d
+ N_XACCXOR/X_XOR8/N002_XACCXOR/X_xor8/M3_g N_GND_XACCXOR/X_xor8/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor10/M3 N_CACC[10]_XACCXOR/X_xor10/M3_d
+ N_XACCXOR/X_XOR10/N002_XACCXOR/X_xor10/M3_g N_GND_XACCXOR/X_xor10/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa72/M2 N_XADDER/XA72/N002_XADDER/Xa72/M2_d
+ N_XADDER/GG1_XADDER/Xa72/M2_g N_XADDER/P2_XADDER/Xa72/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa70/M3 N_OUT1[0]_XADDER/Xa70/M3_d N_XADDER/XA70/N002_XADDER/Xa70/M3_g
+ N_GND_XADDER/Xa70/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa000/Xao2/M37 N_XADDER/XA000/XAO2/N008_XADDER/Xa000/Xao2/M37_d
+ N_XADDER/XA000/OUT1_XADDER/Xa000/Xao2/M37_g N_GND_XADDER/Xa000/Xao2/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xdffa4/M8 N_XBOOTH/XDFFA4/N3_XBOOTH/Xdffa4/M8_d N_CLK_XBOOTH/Xdffa4/M8_g
+ N_XBOOTH/XDFFA4/P003_XBOOTH/Xdffa4/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xdffa5/M8 N_XBOOTH/XDFFA5/N3_XBOOTH/Xdffa5/M8_d N_CLK_XBOOTH/Xdffa5/M8_g
+ N_XBOOTH/XDFFA5/P003_XBOOTH/Xdffa5/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xdffa3/M8 N_XBOOTH/XDFFA3/N3_XBOOTH/Xdffa3/M8_d N_CLK_XBOOTH/Xdffa3/M8_g
+ N_XBOOTH/XDFFA3/P003_XBOOTH/Xdffa3/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xdffa2/M8 N_XBOOTH/XDFFA2/N3_XBOOTH/Xdffa2/M8_d N_CLK_XBOOTH/Xdffa2/M8_g
+ N_XBOOTH/XDFFA2/P003_XBOOTH/Xdffa2/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xdffa0/M8 N_XBOOTH/XDFFA0/N3_XBOOTH/Xdffa0/M8_d N_CLK_XBOOTH/Xdffa0/M8_g
+ N_XBOOTH/XDFFA0/P003_XBOOTH/Xdffa0/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xdffa1/M8 N_XBOOTH/XDFFA1/N3_XBOOTH/Xdffa1/M8_d N_CLK_XBOOTH/Xdffa1/M8_g
+ N_XBOOTH/XDFFA1/P003_XBOOTH/Xdffa1/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa01/Xrb1/M10 N_XADDER/XA01/XRB1/N004_XADDER/Xa01/Xrb1/M10_d
+ N_S[0]_XADDER/Xa01/Xrb1/M10_g N_GND_XADDER/Xa01/Xrb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXACCXOR/X_xor1/M1 N_XACCXOR/X_XOR1/N002_XACCXOR/X_xor1/M1_d
+ N_XACCXOR/DACC[1]_XACCXOR/X_xor1/M1_g N_DMODE_XACCXOR/X_xor1/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXACCXOR/X_xor2/M1 N_XACCXOR/X_XOR2/N002_XACCXOR/X_xor2/M1_d
+ N_XACCXOR/DACC[2]_XACCXOR/X_xor2/M1_g N_DMODE_XACCXOR/X_xor2/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXACCXOR/X_xor4/M1 N_XACCXOR/X_XOR4/N002_XACCXOR/X_xor4/M1_d
+ N_XACCXOR/DACC[4]_XACCXOR/X_xor4/M1_g N_DMODE_XACCXOR/X_xor4/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXACCXOR/X_xor6/M1 N_XACCXOR/X_XOR6/N002_XACCXOR/X_xor6/M1_d
+ N_XACCXOR/DACC[6]_XACCXOR/X_xor6/M1_g N_DMODE_XACCXOR/X_xor6/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXACCXOR/X_xor8/M1 N_XACCXOR/X_XOR8/N002_XACCXOR/X_xor8/M1_d
+ N_XACCXOR/DACC[8]_XACCXOR/X_xor8/M1_g N_DMODE_XACCXOR/X_xor8/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXACCXOR/X_xor10/M1 N_XACCXOR/X_XOR10/N002_XACCXOR/X_xor10/M1_d
+ N_XACCXOR/DACC[10]_XACCXOR/X_xor10/M1_g N_DMODE_XACCXOR/X_xor10/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xdffa4/M9 N_XBOOTH/XDFFA4/P003_XBOOTH/Xdffa4/M9_d
+ N_XBOOTH/XDFFA4/N1_XBOOTH/Xdffa4/M9_g N_GND_XBOOTH/Xdffa4/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXBOOTH/Xdffa5/M9 N_XBOOTH/XDFFA5/P003_XBOOTH/Xdffa5/M9_d
+ N_XBOOTH/XDFFA5/N1_XBOOTH/Xdffa5/M9_g N_GND_XBOOTH/Xdffa5/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXBOOTH/Xdffa3/M9 N_XBOOTH/XDFFA3/P003_XBOOTH/Xdffa3/M9_d
+ N_XBOOTH/XDFFA3/N1_XBOOTH/Xdffa3/M9_g N_GND_XBOOTH/Xdffa3/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXBOOTH/Xdffa2/M9 N_XBOOTH/XDFFA2/P003_XBOOTH/Xdffa2/M9_d
+ N_XBOOTH/XDFFA2/N1_XBOOTH/Xdffa2/M9_g N_GND_XBOOTH/Xdffa2/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXBOOTH/Xdffa0/M9 N_XBOOTH/XDFFA0/P003_XBOOTH/Xdffa0/M9_d
+ N_XBOOTH/XDFFA0/N1_XBOOTH/Xdffa0/M9_g N_GND_XBOOTH/Xdffa0/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXBOOTH/Xdffa1/M9 N_XBOOTH/XDFFA1/P003_XBOOTH/Xdffa1/M9_d
+ N_XBOOTH/XDFFA1/N1_XBOOTH/Xdffa1/M9_g N_GND_XBOOTH/Xdffa1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXADDER/Xa000/Xao2/M38 N_XADDER/XA000/XAO2/N008_XADDER/Xa000/Xao2/M38_d
+ N_XADDER/G0_XADDER/Xa000/Xao2/M38_g N_GND_XADDER/Xa000/Xao2/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa01/Xrb1/M9 N_XADDER/XA01/XRB1/N003_XADDER/Xa01/Xrb1/M9_d
+ N_GND_XADDER/Xa01/Xrb1/M9_g N_XADDER/XA01/XRB1/N004_XADDER/Xa01/Xrb1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14
+ PD=1.44e-06 PS=2.8e-07
mXACCXOR/X_xor1/M2 N_XACCXOR/X_XOR1/N002_XACCXOR/X_xor1/M2_d
+ N_DMODE_XACCXOR/X_xor1/M2_g N_XACCXOR/DACC[1]_XACCXOR/X_xor1/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXACCXOR/X_xor2/M2 N_XACCXOR/X_XOR2/N002_XACCXOR/X_xor2/M2_d
+ N_DMODE_XACCXOR/X_xor2/M2_g N_XACCXOR/DACC[2]_XACCXOR/X_xor2/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXACCXOR/X_xor4/M2 N_XACCXOR/X_XOR4/N002_XACCXOR/X_xor4/M2_d
+ N_DMODE_XACCXOR/X_xor4/M2_g N_XACCXOR/DACC[4]_XACCXOR/X_xor4/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXACCXOR/X_xor6/M2 N_XACCXOR/X_XOR6/N002_XACCXOR/X_xor6/M2_d
+ N_DMODE_XACCXOR/X_xor6/M2_g N_XACCXOR/DACC[6]_XACCXOR/X_xor6/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXACCXOR/X_xor8/M2 N_XACCXOR/X_XOR8/N002_XACCXOR/X_xor8/M2_d
+ N_DMODE_XACCXOR/X_xor8/M2_g N_XACCXOR/DACC[8]_XACCXOR/X_xor8/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXACCXOR/X_xor10/M2 N_XACCXOR/X_XOR10/N002_XACCXOR/X_xor10/M2_d
+ N_DMODE_XACCXOR/X_xor10/M2_g N_XACCXOR/DACC[10]_XACCXOR/X_xor10/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mX02/xd21/M3 N_X02/XD21/N0_X02/xd21/M3_d N_OUT1[0]_X02/xd21/M3_g
+ N_GND_X02/xd21/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXADDER/Xa73/M3 N_OUT1[3]_XADDER/Xa73/M3_d N_XADDER/XA73/N002_XADDER/Xa73/M3_g
+ N_GND_XADDER/Xa73/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xdffa4/M11 N_XBOOTH/A_D[4]_XBOOTH/Xdffa4/M11_d
+ N_XBOOTH/XDFFA4/N3_XBOOTH/Xdffa4/M11_g N_GND_XBOOTH/Xdffa4/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXBOOTH/Xdffa5/M11 N_A_D[5]_XBOOTH/Xdffa5/M11_d
+ N_XBOOTH/XDFFA5/N3_XBOOTH/Xdffa5/M11_g N_GND_XBOOTH/Xdffa5/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXBOOTH/Xdffa3/M11 N_A_D[3]_XBOOTH/Xdffa3/M11_d
+ N_XBOOTH/XDFFA3/N3_XBOOTH/Xdffa3/M11_g N_GND_XBOOTH/Xdffa3/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXBOOTH/Xdffa2/M11 N_XBOOTH/A_D[2]_XBOOTH/Xdffa2/M11_d
+ N_XBOOTH/XDFFA2/N3_XBOOTH/Xdffa2/M11_g N_GND_XBOOTH/Xdffa2/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXBOOTH/Xdffa0/M11 N_XBOOTH/A_D[0]_XBOOTH/Xdffa0/M11_d
+ N_XBOOTH/XDFFA0/N3_XBOOTH/Xdffa0/M11_g N_GND_XBOOTH/Xdffa0/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXBOOTH/Xdffa1/M11 N_A_D[1]_XBOOTH/Xdffa1/M11_d
+ N_XBOOTH/XDFFA1/N3_XBOOTH/Xdffa1/M11_g N_GND_XBOOTH/Xdffa1/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mX02/xd21/M6 N_X02/XD21/P002_X02/xd21/M6_d N_CLK_X02/xd21/M6_g
+ N_GND_X02/xd21/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXADDER/Xa000/Xao2/Xor1/M16 N_XADDER/G00_XADDER/Xa000/Xao2/Xor1/M16_d
+ N_XADDER/XA000/XAO2/N008_XADDER/Xa000/Xao2/Xor1/M16_g
+ N_GND_XADDER/Xa000/Xao2/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa01/Xrb1/Xand1/M16 N_XADDER/G0_XADDER/Xa01/Xrb1/Xand1/M16_d
+ N_XADDER/XA01/XRB1/N003_XADDER/Xa01/Xrb1/Xand1/M16_g
+ N_GND_XADDER/Xa01/Xrb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd21/M5 N_X02/XD21/N1_X02/xd21/M5_d N_X02/XD21/N0_X02/xd21/M5_g
+ N_X02/XD21/P002_X02/xd21/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa12/M3 N_XACCXOR/XDFFA12/N0_XACCXOR/Xdffa12/M3_d
+ N_MODE_XACCXOR/Xdffa12/M3_g N_GND_XACCXOR/Xdffa12/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa71/M2 N_XADDER/XA71/N002_XADDER/Xa71/M2_d
+ N_XADDER/G00_XADDER/Xa71/M2_g N_XADDER/P1_XADDER/Xa71/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXACCXOR/Xdffa1/M11 N_XACCXOR/DACC[1]_XACCXOR/Xdffa1/M11_d
+ N_XACCXOR/XDFFA1/N3_XACCXOR/Xdffa1/M11_g N_GND_XACCXOR/Xdffa1/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXACCXOR/Xdffa2/M11 N_XACCXOR/DACC[2]_XACCXOR/Xdffa2/M11_d
+ N_XACCXOR/XDFFA2/N3_XACCXOR/Xdffa2/M11_g N_GND_XACCXOR/Xdffa2/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXACCXOR/Xdffa4/M11 N_XACCXOR/DACC[4]_XACCXOR/Xdffa4/M11_d
+ N_XACCXOR/XDFFA4/N3_XACCXOR/Xdffa4/M11_g N_GND_XACCXOR/Xdffa4/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXACCXOR/Xdffa6/M11 N_XACCXOR/DACC[6]_XACCXOR/Xdffa6/M11_d
+ N_XACCXOR/XDFFA6/N3_XACCXOR/Xdffa6/M11_g N_GND_XACCXOR/Xdffa6/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXACCXOR/Xdffa8/M11 N_XACCXOR/DACC[8]_XACCXOR/Xdffa8/M11_d
+ N_XACCXOR/XDFFA8/N3_XACCXOR/Xdffa8/M11_g N_GND_XACCXOR/Xdffa8/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXACCXOR/Xdffa10/M11 N_XACCXOR/DACC[10]_XACCXOR/Xdffa10/M11_d
+ N_XACCXOR/XDFFA10/N3_XACCXOR/Xdffa10/M11_g N_GND_XACCXOR/Xdffa10/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXACCXOR/Xdffa12/M6 N_XACCXOR/XDFFA12/P002_XACCXOR/Xdffa12/M6_d
+ N_CLK_XACCXOR/Xdffa12/M6_g N_GND_XACCXOR/Xdffa12/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXADDER/Xa71/M1 N_XADDER/XA71/N002_XADDER/Xa71/M1_d N_XADDER/P1_XADDER/Xa71/M1_g
+ N_XADDER/G00_XADDER/Xa71/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=2.332e-13 PD=5.4e-07 PS=1.5e-06
mXADDER/Xa73/M1 N_XADDER/XA73/N002_XADDER/Xa73/M1_d N_XADDER/P3_XADDER/Xa73/M1_g
+ N_XADDER/GX6[0]_XADDER/Xa73/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=2.332e-13 PD=5.4e-07 PS=1.5e-06
mXBOOTH/Xe2/M8 N_XBOOTH/XE2/_B_XBOOTH/Xe2/M8_d N_XBOOTH/A_D[4]_XBOOTH/Xe2/M8_g
+ N_GND_XBOOTH/Xe2/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe1/M8 N_XBOOTH/XE1/_B_XBOOTH/Xe1/M8_d N_XBOOTH/A_D[2]_XBOOTH/Xe1/M8_g
+ N_GND_XBOOTH/Xe1/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe0/M8 N_XBOOTH/XE0/_B_XBOOTH/Xe0/M8_d N_XBOOTH/A_D[0]_XBOOTH/Xe0/M8_g
+ N_GND_XBOOTH/Xe0/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa12/M5 N_XACCXOR/XDFFA12/N1_XACCXOR/Xdffa12/M5_d
+ N_XACCXOR/XDFFA12/N0_XACCXOR/Xdffa12/M5_g
+ N_XACCXOR/XDFFA12/P002_XACCXOR/Xdffa12/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa1/M9 N_XACCXOR/XDFFA1/P003_XACCXOR/Xdffa1/M9_d
+ N_XACCXOR/XDFFA1/N1_XACCXOR/Xdffa1/M9_g N_GND_XACCXOR/Xdffa1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXACCXOR/Xdffa2/M9 N_XACCXOR/XDFFA2/P003_XACCXOR/Xdffa2/M9_d
+ N_XACCXOR/XDFFA2/N1_XACCXOR/Xdffa2/M9_g N_GND_XACCXOR/Xdffa2/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXACCXOR/Xdffa4/M9 N_XACCXOR/XDFFA4/P003_XACCXOR/Xdffa4/M9_d
+ N_XACCXOR/XDFFA4/N1_XACCXOR/Xdffa4/M9_g N_GND_XACCXOR/Xdffa4/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXACCXOR/Xdffa6/M9 N_XACCXOR/XDFFA6/P003_XACCXOR/Xdffa6/M9_d
+ N_XACCXOR/XDFFA6/N1_XACCXOR/Xdffa6/M9_g N_GND_XACCXOR/Xdffa6/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXACCXOR/Xdffa8/M9 N_XACCXOR/XDFFA8/P003_XACCXOR/Xdffa8/M9_d
+ N_XACCXOR/XDFFA8/N1_XACCXOR/Xdffa8/M9_g N_GND_XACCXOR/Xdffa8/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXACCXOR/Xdffa10/M9 N_XACCXOR/XDFFA10/P003_XACCXOR/Xdffa10/M9_d
+ N_XACCXOR/XDFFA10/N1_XACCXOR/Xdffa10/M9_g N_GND_XACCXOR/Xdffa10/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXADDER/Xa02/Xrb2/M3 N_XADDER/P1_XADDER/Xa02/Xrb2/M3_d
+ N_XADDER/XA02/XRB2/N002_XADDER/Xa02/Xrb2/M3_g N_GND_XADDER/Xa02/Xrb2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa11/Xyb1/Xand1/M16 N_XADDER/PP1_XADDER/Xa11/Xyb1/Xand1/M16_d
+ N_XADDER/XA11/XYB1/N003_XADDER/Xa11/Xyb1/Xand1/M16_g
+ N_GND_XADDER/Xa11/Xyb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd21/M8 N_X02/XD21/N3_X02/xd21/M8_d N_CLK_X02/xd21/M8_g
+ N_X02/XD21/P003_X02/xd21/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa73/M2 N_XADDER/XA73/N002_XADDER/Xa73/M2_d
+ N_XADDER/GX6[0]_XADDER/Xa73/M2_g N_XADDER/P3_XADDER/Xa73/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXACCXOR/Xdffa1/M8 N_XACCXOR/XDFFA1/N3_XACCXOR/Xdffa1/M8_d
+ N_CLK_XACCXOR/Xdffa1/M8_g N_XACCXOR/XDFFA1/P003_XACCXOR/Xdffa1/M8_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa2/M8 N_XACCXOR/XDFFA2/N3_XACCXOR/Xdffa2/M8_d
+ N_CLK_XACCXOR/Xdffa2/M8_g N_XACCXOR/XDFFA2/P003_XACCXOR/Xdffa2/M8_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa4/M8 N_XACCXOR/XDFFA4/N3_XACCXOR/Xdffa4/M8_d
+ N_CLK_XACCXOR/Xdffa4/M8_g N_XACCXOR/XDFFA4/P003_XACCXOR/Xdffa4/M8_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa6/M8 N_XACCXOR/XDFFA6/N3_XACCXOR/Xdffa6/M8_d
+ N_CLK_XACCXOR/Xdffa6/M8_g N_XACCXOR/XDFFA6/P003_XACCXOR/Xdffa6/M8_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa8/M8 N_XACCXOR/XDFFA8/N3_XACCXOR/Xdffa8/M8_d
+ N_CLK_XACCXOR/Xdffa8/M8_g N_XACCXOR/XDFFA8/P003_XACCXOR/Xdffa8/M8_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa10/M8 N_XACCXOR/XDFFA10/N3_XACCXOR/Xdffa10/M8_d
+ N_CLK_XACCXOR/Xdffa10/M8_g N_XACCXOR/XDFFA10/P003_XACCXOR/Xdffa10/M8_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xe2/M7 N_XBOOTH/XE2/_A_XBOOTH/Xe2/M7_d N_A_D[5]_XBOOTH/Xe2/M7_g
+ N_GND_XBOOTH/Xe2/M7_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.464e-13 AS=1.188e-13 PD=1.56e-06 PS=5.4e-07
mXBOOTH/Xe1/M7 N_XBOOTH/XE1/_A_XBOOTH/Xe1/M7_d N_A_D[3]_XBOOTH/Xe1/M7_g
+ N_GND_XBOOTH/Xe1/M7_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.464e-13 AS=1.188e-13 PD=1.56e-06 PS=5.4e-07
mXBOOTH/Xe0/M7 N_XBOOTH/XE0/_A_XBOOTH/Xe0/M7_d N_A_D[1]_XBOOTH/Xe0/M7_g
+ N_GND_XBOOTH/Xe0/M7_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.464e-13 AS=1.188e-13 PD=1.56e-06 PS=5.4e-07
mX02/xd21/M9 N_X02/XD21/P003_X02/xd21/M9_d N_X02/XD21/N1_X02/xd21/M9_g
+ N_GND_X02/xd21/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.76e-13 PD=2.8e-07 PS=8e-07
mXACCXOR/Xdffa12/M8 N_XACCXOR/XDFFA12/N3_XACCXOR/Xdffa12/M8_d
+ N_CLK_XACCXOR/Xdffa12/M8_g N_XACCXOR/XDFFA12/P003_XACCXOR/Xdffa12/M8_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa71/M3 N_OUT1[1]_XADDER/Xa71/M3_d N_XADDER/XA71/N002_XADDER/Xa71/M3_g
+ N_GND_XADDER/Xa71/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa02/Xrb2/M1 N_XADDER/XA02/XRB2/N002_XADDER/Xa02/Xrb2/M1_d
+ N_C[1]_XADDER/Xa02/Xrb2/M1_g N_S[1]_XADDER/Xa02/Xrb2/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa11/Xyb1/M9 N_XADDER/XA11/XYB1/N003_XADDER/Xa11/Xyb1/M9_d
+ N_XADDER/P0_XADDER/Xa11/Xyb1/M9_g
+ N_XADDER/XA11/XYB1/N004_XADDER/Xa11/Xyb1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=9.24e-14 PD=1.44e-06 PS=4.2e-07
mX02/xd21/M11 N_OUT[0]_X02/xd21/M11_d N_X02/XD21/N3_X02/xd21/M11_g
+ N_GND_X02/xd21/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXACCXOR/Xdffa12/M9 N_XACCXOR/XDFFA12/P003_XACCXOR/Xdffa12/M9_d
+ N_XACCXOR/XDFFA12/N1_XACCXOR/Xdffa12/M9_g N_GND_XACCXOR/Xdffa12/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXACCXOR/Xdffa1/M5 N_XACCXOR/XDFFA1/N1_XACCXOR/Xdffa1/M5_d
+ N_XACCXOR/XDFFA1/N0_XACCXOR/Xdffa1/M5_g
+ N_XACCXOR/XDFFA1/P002_XACCXOR/Xdffa1/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa2/M5 N_XACCXOR/XDFFA2/N1_XACCXOR/Xdffa2/M5_d
+ N_XACCXOR/XDFFA2/N0_XACCXOR/Xdffa2/M5_g
+ N_XACCXOR/XDFFA2/P002_XACCXOR/Xdffa2/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa4/M5 N_XACCXOR/XDFFA4/N1_XACCXOR/Xdffa4/M5_d
+ N_XACCXOR/XDFFA4/N0_XACCXOR/Xdffa4/M5_g
+ N_XACCXOR/XDFFA4/P002_XACCXOR/Xdffa4/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa6/M5 N_XACCXOR/XDFFA6/N1_XACCXOR/Xdffa6/M5_d
+ N_XACCXOR/XDFFA6/N0_XACCXOR/Xdffa6/M5_g
+ N_XACCXOR/XDFFA6/P002_XACCXOR/Xdffa6/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa8/M5 N_XACCXOR/XDFFA8/N1_XACCXOR/Xdffa8/M5_d
+ N_XACCXOR/XDFFA8/N0_XACCXOR/Xdffa8/M5_g
+ N_XACCXOR/XDFFA8/P002_XACCXOR/Xdffa8/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa10/M5 N_XACCXOR/XDFFA10/N1_XACCXOR/Xdffa10/M5_d
+ N_XACCXOR/XDFFA10/N0_XACCXOR/Xdffa10/M5_g
+ N_XACCXOR/XDFFA10/P002_XACCXOR/Xdffa10/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xe2/M6 N_noxref_2070_XBOOTH/Xe2/M6_d N_A_D[5]_XBOOTH/Xe2/M6_g
+ N_GND_XBOOTH/Xe2/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xe2/M1 N_noxref_2071_XBOOTH/Xe2/M1_d N_XBOOTH/XE2/_A_XBOOTH/Xe2/M1_g
+ N_GND_XBOOTH/Xe2/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xe1/M1 N_noxref_2072_XBOOTH/Xe1/M1_d N_XBOOTH/XE1/_A_XBOOTH/Xe1/M1_g
+ N_GND_XBOOTH/Xe1/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xe1/M6 N_noxref_2073_XBOOTH/Xe1/M6_d N_A_D[3]_XBOOTH/Xe1/M6_g
+ N_GND_XBOOTH/Xe1/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xe0/M6 N_noxref_2074_XBOOTH/Xe0/M6_d N_A_D[1]_XBOOTH/Xe0/M6_g
+ N_GND_XBOOTH/Xe0/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xe0/M1 N_noxref_2075_XBOOTH/Xe0/M1_d N_XBOOTH/XE0/_A_XBOOTH/Xe0/M1_g
+ N_GND_XBOOTH/Xe0/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXADDER/Xa74/M3 N_OUT1[4]_XADDER/Xa74/M3_d N_XADDER/XA74/N002_XADDER/Xa74/M3_g
+ N_GND_XADDER/Xa74/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa11/Xyb1/M10 N_XADDER/XA11/XYB1/N004_XADDER/Xa11/Xyb1/M10_d
+ N_XADDER/P1_XADDER/Xa11/Xyb1/M10_g N_GND_XADDER/Xa11/Xyb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=9.24e-14 AS=2.244e-13
+ PD=4.2e-07 PS=1.46e-06
mXADDER/Xa02/Xrb2/M2 N_XADDER/XA02/XRB2/N002_XADDER/Xa02/Xrb2/M2_d
+ N_S[1]_XADDER/Xa02/Xrb2/M2_g N_C[1]_XADDER/Xa02/Xrb2/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXACCXOR/Xdffa1/M6 N_XACCXOR/XDFFA1/P002_XACCXOR/Xdffa1/M6_d
+ N_CLK_XACCXOR/Xdffa1/M6_g N_GND_XACCXOR/Xdffa1/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXACCXOR/Xdffa2/M6 N_XACCXOR/XDFFA2/P002_XACCXOR/Xdffa2/M6_d
+ N_CLK_XACCXOR/Xdffa2/M6_g N_GND_XACCXOR/Xdffa2/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXACCXOR/Xdffa4/M6 N_XACCXOR/XDFFA4/P002_XACCXOR/Xdffa4/M6_d
+ N_CLK_XACCXOR/Xdffa4/M6_g N_GND_XACCXOR/Xdffa4/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXACCXOR/Xdffa6/M6 N_XACCXOR/XDFFA6/P002_XACCXOR/Xdffa6/M6_d
+ N_CLK_XACCXOR/Xdffa6/M6_g N_GND_XACCXOR/Xdffa6/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXACCXOR/Xdffa8/M6 N_XACCXOR/XDFFA8/P002_XACCXOR/Xdffa8/M6_d
+ N_CLK_XACCXOR/Xdffa8/M6_g N_GND_XACCXOR/Xdffa8/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXACCXOR/Xdffa10/M6 N_XACCXOR/XDFFA10/P002_XACCXOR/Xdffa10/M6_d
+ N_CLK_XACCXOR/Xdffa10/M6_g N_GND_XACCXOR/Xdffa10/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXBOOTH/Xe2/M5 N_noxref_2076_XBOOTH/Xe2/M5_d N_XBOOTH/XE2/_B_XBOOTH/Xe2/M5_g
+ N_noxref_2070_XBOOTH/Xe2/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=1.188e-13 PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xe2/M2 N_noxref_2077_XBOOTH/Xe2/M2_d N_XBOOTH/A_D[4]_XBOOTH/Xe2/M2_g
+ N_noxref_2071_XBOOTH/Xe2/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=1.188e-13 PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xe1/M2 N_noxref_2078_XBOOTH/Xe1/M2_d N_XBOOTH/A_D[2]_XBOOTH/Xe1/M2_g
+ N_noxref_2072_XBOOTH/Xe1/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=1.188e-13 PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xe1/M5 N_noxref_2079_XBOOTH/Xe1/M5_d N_XBOOTH/XE1/_B_XBOOTH/Xe1/M5_g
+ N_noxref_2073_XBOOTH/Xe1/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=1.188e-13 PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xe0/M5 N_noxref_2080_XBOOTH/Xe0/M5_d N_XBOOTH/XE0/_B_XBOOTH/Xe0/M5_g
+ N_noxref_2074_XBOOTH/Xe0/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=1.188e-13 PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xe0/M2 N_noxref_2081_XBOOTH/Xe0/M2_d N_XBOOTH/A_D[0]_XBOOTH/Xe0/M2_g
+ N_noxref_2075_XBOOTH/Xe0/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=1.188e-13 PD=5.4e-07 PS=5.4e-07
mXACCXOR/Xdffa12/M11 N_DMODE_XACCXOR/Xdffa12/M11_d
+ N_XACCXOR/XDFFA12/N3_XACCXOR/Xdffa12/M11_g N_GND_XACCXOR/Xdffa12/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mX02/xd22/M3 N_X02/XD22/N0_X02/xd22/M3_d N_OUT1[1]_X02/xd22/M3_g
+ N_GND_X02/xd22/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXADDER/Xa62/Xao2/Xor1/M16 N_XADDER/GX6[0]_XADDER/Xa62/Xao2/Xor1/M16_d
+ N_XADDER/XA62/XAO2/N008_XADDER/Xa62/Xao2/Xor1/M16_g
+ N_GND_XADDER/Xa62/Xao2/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXACCXOR/Xdffa1/M3 N_XACCXOR/XDFFA1/N0_XACCXOR/Xdffa1/M3_d
+ N_ACC[1]_XACCXOR/Xdffa1/M3_g N_GND_XACCXOR/Xdffa1/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa2/M3 N_XACCXOR/XDFFA2/N0_XACCXOR/Xdffa2/M3_d
+ N_ACC[2]_XACCXOR/Xdffa2/M3_g N_GND_XACCXOR/Xdffa2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa4/M3 N_XACCXOR/XDFFA4/N0_XACCXOR/Xdffa4/M3_d
+ N_ACC[4]_XACCXOR/Xdffa4/M3_g N_GND_XACCXOR/Xdffa4/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa6/M3 N_XACCXOR/XDFFA6/N0_XACCXOR/Xdffa6/M3_d
+ N_ACC[6]_XACCXOR/Xdffa6/M3_g N_GND_XACCXOR/Xdffa6/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa8/M3 N_XACCXOR/XDFFA8/N0_XACCXOR/Xdffa8/M3_d
+ N_ACC[8]_XACCXOR/Xdffa8/M3_g N_GND_XACCXOR/Xdffa8/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa10/M3 N_XACCXOR/XDFFA10/N0_XACCXOR/Xdffa10/M3_d
+ N_ACC[10]_XACCXOR/Xdffa10/M3_g N_GND_XACCXOR/Xdffa10/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe2/M4 N_XBOOTH/XE2/N002_XBOOTH/Xe2/M4_d N_XBOOTH/XE2/_C_XBOOTH/Xe2/M4_g
+ N_noxref_2076_XBOOTH/Xe2/M4_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe2/M3 N_XBOOTH/XE2/N002_XBOOTH/Xe2/M3_d N_A_D[3]_XBOOTH/Xe2/M3_g
+ N_noxref_2077_XBOOTH/Xe2/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe1/M3 N_XBOOTH/XE1/N002_XBOOTH/Xe1/M3_d N_A_D[1]_XBOOTH/Xe1/M3_g
+ N_noxref_2078_XBOOTH/Xe1/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe1/M4 N_XBOOTH/XE1/N002_XBOOTH/Xe1/M4_d N_XBOOTH/XE1/_C_XBOOTH/Xe1/M4_g
+ N_noxref_2079_XBOOTH/Xe1/M4_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe0/M4 N_XBOOTH/XE0/N002_XBOOTH/Xe0/M4_d N_XBOOTH/XE0/_C_XBOOTH/Xe0/M4_g
+ N_noxref_2080_XBOOTH/Xe0/M4_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe0/M3 N_XBOOTH/XE0/N002_XBOOTH/Xe0/M3_d N_GND_XBOOTH/Xe0/M3_g
+ N_noxref_2081_XBOOTH/Xe0/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXADDER/Xa11/Xyb2/M10 N_XADDER/XA11/XYB2/N004_XADDER/Xa11/Xyb2/M10_d
+ N_XADDER/P1_XADDER/Xa11/Xyb2/M10_g N_GND_XADDER/Xa11/Xyb2/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mX02/xd22/M6 N_X02/XD22/P002_X02/xd22/M6_d N_CLK_X02/xd22/M6_g
+ N_GND_X02/xd22/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXADDER/Xa02/Xrb1/M10 N_XADDER/XA02/XRB1/N004_XADDER/Xa02/Xrb1/M10_d
+ N_S[1]_XADDER/Xa02/Xrb1/M10_g N_GND_XADDER/Xa02/Xrb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXADDER/Xa74/M1 N_XADDER/XA74/N002_XADDER/Xa74/M1_d N_XADDER/P4_XADDER/Xa74/M1_g
+ N_XADDER/GGG3_XADDER/Xa74/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=2.332e-13 PD=5.4e-07 PS=1.5e-06
mXADDER/Xa11/Xyb2/M9 N_XADDER/XA11/XYB2/N003_XADDER/Xa11/Xyb2/M9_d
+ N_XADDER/G00_XADDER/Xa11/Xyb2/M9_g
+ N_XADDER/XA11/XYB2/N004_XADDER/Xa11/Xyb2/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=6.16e-14 PD=1.74e-06 PS=2.8e-07
mX02/xd22/M5 N_X02/XD22/N1_X02/xd22/M5_d N_X02/XD22/N0_X02/xd22/M5_g
+ N_X02/XD22/P002_X02/xd22/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa02/Xrb1/M9 N_XADDER/XA02/XRB1/N003_XADDER/Xa02/Xrb1/M9_d
+ N_C[1]_XADDER/Xa02/Xrb1/M9_g N_XADDER/XA02/XRB1/N004_XADDER/Xa02/Xrb1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14
+ PD=1.44e-06 PS=2.8e-07
mXADDER/Xa62/Xao2/M38 N_XADDER/XA62/XAO2/N008_XADDER/Xa62/Xao2/M38_d
+ N_XADDER/G2_XADDER/Xa62/Xao2/M38_g N_GND_XADDER/Xa62/Xao2/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa0/M3 N_XACCXOR/XDFFA0/N0_XACCXOR/Xdffa0/M3_d
+ N_ACC[0]_XACCXOR/Xdffa0/M3_g N_GND_XACCXOR/Xdffa0/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa3/M3 N_XACCXOR/XDFFA3/N0_XACCXOR/Xdffa3/M3_d
+ N_ACC[3]_XACCXOR/Xdffa3/M3_g N_GND_XACCXOR/Xdffa3/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa5/M3 N_XACCXOR/XDFFA5/N0_XACCXOR/Xdffa5/M3_d
+ N_ACC[5]_XACCXOR/Xdffa5/M3_g N_GND_XACCXOR/Xdffa5/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa7/M3 N_XACCXOR/XDFFA7/N0_XACCXOR/Xdffa7/M3_d
+ N_ACC[7]_XACCXOR/Xdffa7/M3_g N_GND_XACCXOR/Xdffa7/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa9/M3 N_XACCXOR/XDFFA9/N0_XACCXOR/Xdffa9/M3_d
+ N_ACC[9]_XACCXOR/Xdffa9/M3_g N_GND_XACCXOR/Xdffa9/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa11/M3 N_XACCXOR/XDFFA11/N0_XACCXOR/Xdffa11/M3_d
+ N_ACC[11]_XACCXOR/Xdffa11/M3_g N_GND_XACCXOR/Xdffa11/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa74/M2 N_XADDER/XA74/N002_XADDER/Xa74/M2_d
+ N_XADDER/GGG3_XADDER/Xa74/M2_g N_XADDER/P4_XADDER/Xa74/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xe2/M9 N_XBOOTH/XE2/_C_XBOOTH/Xe2/M9_d N_A_D[3]_XBOOTH/Xe2/M9_g
+ N_GND_XBOOTH/Xe2/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.298e-13 PD=1.42e-06 PS=5.9e-07
mXBOOTH/Xe1/M9 N_XBOOTH/XE1/_C_XBOOTH/Xe1/M9_d N_A_D[1]_XBOOTH/Xe1/M9_g
+ N_GND_XBOOTH/Xe1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.298e-13 PD=1.42e-06 PS=5.9e-07
mXBOOTH/Xe0/M9 N_XBOOTH/XE0/_C_XBOOTH/Xe0/M9_d N_GND_XBOOTH/Xe0/M9_g
+ N_GND_XBOOTH/Xe0/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.298e-13 PD=1.42e-06 PS=5.9e-07
mXADDER/Xa62/Xao2/M37 N_XADDER/XA62/XAO2/N008_XADDER/Xa62/Xao2/M37_d
+ N_XADDER/XA62/OUT1_XADDER/Xa62/Xao2/M37_g N_GND_XADDER/Xa62/Xao2/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa0/M6 N_XACCXOR/XDFFA0/P002_XACCXOR/Xdffa0/M6_d
+ N_CLK_XACCXOR/Xdffa0/M6_g N_GND_XACCXOR/Xdffa0/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXACCXOR/Xdffa3/M6 N_XACCXOR/XDFFA3/P002_XACCXOR/Xdffa3/M6_d
+ N_CLK_XACCXOR/Xdffa3/M6_g N_GND_XACCXOR/Xdffa3/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXACCXOR/Xdffa5/M6 N_XACCXOR/XDFFA5/P002_XACCXOR/Xdffa5/M6_d
+ N_CLK_XACCXOR/Xdffa5/M6_g N_GND_XACCXOR/Xdffa5/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXACCXOR/Xdffa7/M6 N_XACCXOR/XDFFA7/P002_XACCXOR/Xdffa7/M6_d
+ N_CLK_XACCXOR/Xdffa7/M6_g N_GND_XACCXOR/Xdffa7/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXACCXOR/Xdffa9/M6 N_XACCXOR/XDFFA9/P002_XACCXOR/Xdffa9/M6_d
+ N_CLK_XACCXOR/Xdffa9/M6_g N_GND_XACCXOR/Xdffa9/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXACCXOR/Xdffa11/M6 N_XACCXOR/XDFFA11/P002_XACCXOR/Xdffa11/M6_d
+ N_CLK_XACCXOR/Xdffa11/M6_g N_GND_XACCXOR/Xdffa11/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mX02/xd22/M8 N_X02/XD22/N3_X02/xd22/M8_d N_CLK_X02/xd22/M8_g
+ N_X02/XD22/P003_X02/xd22/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa0/M5 N_XACCXOR/XDFFA0/N1_XACCXOR/Xdffa0/M5_d
+ N_XACCXOR/XDFFA0/N0_XACCXOR/Xdffa0/M5_g
+ N_XACCXOR/XDFFA0/P002_XACCXOR/Xdffa0/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa3/M5 N_XACCXOR/XDFFA3/N1_XACCXOR/Xdffa3/M5_d
+ N_XACCXOR/XDFFA3/N0_XACCXOR/Xdffa3/M5_g
+ N_XACCXOR/XDFFA3/P002_XACCXOR/Xdffa3/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa5/M5 N_XACCXOR/XDFFA5/N1_XACCXOR/Xdffa5/M5_d
+ N_XACCXOR/XDFFA5/N0_XACCXOR/Xdffa5/M5_g
+ N_XACCXOR/XDFFA5/P002_XACCXOR/Xdffa5/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa7/M5 N_XACCXOR/XDFFA7/N1_XACCXOR/Xdffa7/M5_d
+ N_XACCXOR/XDFFA7/N0_XACCXOR/Xdffa7/M5_g
+ N_XACCXOR/XDFFA7/P002_XACCXOR/Xdffa7/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa9/M5 N_XACCXOR/XDFFA9/N1_XACCXOR/Xdffa9/M5_d
+ N_XACCXOR/XDFFA9/N0_XACCXOR/Xdffa9/M5_g
+ N_XACCXOR/XDFFA9/P002_XACCXOR/Xdffa9/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa11/M5 N_XACCXOR/XDFFA11/N1_XACCXOR/Xdffa11/M5_d
+ N_XACCXOR/XDFFA11/N0_XACCXOR/Xdffa11/M5_g
+ N_XACCXOR/XDFFA11/P002_XACCXOR/Xdffa11/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa11/Xyb2/Xand1/M16 N_XADDER/XA11/T1_XADDER/Xa11/Xyb2/Xand1/M16_d
+ N_XADDER/XA11/XYB2/N003_XADDER/Xa11/Xyb2/Xand1/M16_g
+ N_GND_XADDER/Xa11/Xyb2/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xe2/M19 N_XBOOTH/D2_XBOOTH/Xe2/M19_d N_XBOOTH/XE2/N002_XBOOTH/Xe2/M19_g
+ N_GND_XBOOTH/Xe2/M19_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.298e-13 PD=1.42e-06 PS=5.9e-07
mXBOOTH/Xe1/M19 N_XBOOTH/D1_XBOOTH/Xe1/M19_d N_XBOOTH/XE1/N002_XBOOTH/Xe1/M19_g
+ N_GND_XBOOTH/Xe1/M19_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.298e-13 PD=1.42e-06 PS=5.9e-07
mXBOOTH/Xe0/M19 N_XBOOTH/D0_XBOOTH/Xe0/M19_d N_XBOOTH/XE0/N002_XBOOTH/Xe0/M19_g
+ N_GND_XBOOTH/Xe0/M19_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.298e-13 PD=1.42e-06 PS=5.9e-07
mXADDER/Xa02/Xrb1/Xand1/M16 N_XADDER/G1_XADDER/Xa02/Xrb1/Xand1/M16_d
+ N_XADDER/XA02/XRB1/N003_XADDER/Xa02/Xrb1/Xand1/M16_g
+ N_GND_XADDER/Xa02/Xrb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd22/M9 N_X02/XD22/P003_X02/xd22/M9_d N_X02/XD22/N1_X02/xd22/M9_g
+ N_GND_X02/xd22/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.76e-13 PD=2.8e-07 PS=8e-07
mXADDER/Xa62/Xao1/Xand1/M16 N_XADDER/XA62/OUT1_XADDER/Xa62/Xao1/Xand1/M16_d
+ N_XADDER/XA62/XAO1/N003_XADDER/Xa62/Xao1/Xand1/M16_g
+ N_GND_XADDER/Xa62/Xao1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd22/M11 N_OUT[1]_X02/xd22/M11_d N_X02/XD22/N3_X02/xd22/M11_g
+ N_GND_X02/xd22/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXACCXOR/Xdffa0/M8 N_XACCXOR/XDFFA0/N3_XACCXOR/Xdffa0/M8_d
+ N_CLK_XACCXOR/Xdffa0/M8_g N_XACCXOR/XDFFA0/P003_XACCXOR/Xdffa0/M8_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa3/M8 N_XACCXOR/XDFFA3/N3_XACCXOR/Xdffa3/M8_d
+ N_CLK_XACCXOR/Xdffa3/M8_g N_XACCXOR/XDFFA3/P003_XACCXOR/Xdffa3/M8_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa5/M8 N_XACCXOR/XDFFA5/N3_XACCXOR/Xdffa5/M8_d
+ N_CLK_XACCXOR/Xdffa5/M8_g N_XACCXOR/XDFFA5/P003_XACCXOR/Xdffa5/M8_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa7/M8 N_XACCXOR/XDFFA7/N3_XACCXOR/Xdffa7/M8_d
+ N_CLK_XACCXOR/Xdffa7/M8_g N_XACCXOR/XDFFA7/P003_XACCXOR/Xdffa7/M8_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa9/M8 N_XACCXOR/XDFFA9/N3_XACCXOR/Xdffa9/M8_d
+ N_CLK_XACCXOR/Xdffa9/M8_g N_XACCXOR/XDFFA9/P003_XACCXOR/Xdffa9/M8_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa11/M8 N_XACCXOR/XDFFA11/N3_XACCXOR/Xdffa11/M8_d
+ N_CLK_XACCXOR/Xdffa11/M8_g N_XACCXOR/XDFFA11/P003_XACCXOR/Xdffa11/M8_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa11/Xyb3/M37 N_XADDER/XA11/XYB3/N008_XADDER/Xa11/Xyb3/M37_d
+ N_XADDER/XA11/T1_XADDER/Xa11/Xyb3/M37_g N_GND_XADDER/Xa11/Xyb3/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe2/M22 N_XBOOTH/XE2/N004_XBOOTH/Xe2/M22_d N_A_D[3]_XBOOTH/Xe2/M22_g
+ N_XBOOTH/A_D[4]_XBOOTH/Xe2/M22_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=2.2e-13 PD=5.4e-07 PS=1.44e-06
mXBOOTH/Xe1/M22 N_XBOOTH/XE1/N004_XBOOTH/Xe1/M22_d N_A_D[1]_XBOOTH/Xe1/M22_g
+ N_XBOOTH/A_D[2]_XBOOTH/Xe1/M22_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=2.2e-13 PD=5.4e-07 PS=1.44e-06
mXBOOTH/Xe0/M22 N_XBOOTH/XE0/N004_XBOOTH/Xe0/M22_d N_GND_XBOOTH/Xe0/M22_g
+ N_XBOOTH/A_D[0]_XBOOTH/Xe0/M22_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=2.2e-13 PD=5.4e-07 PS=1.44e-06
mXADDER/Xa03/Xrb2/M3 N_XADDER/P2_XADDER/Xa03/Xrb2/M3_d
+ N_XADDER/XA03/XRB2/N002_XADDER/Xa03/Xrb2/M3_g N_GND_XADDER/Xa03/Xrb2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/Xdffa0/M9 N_XACCXOR/XDFFA0/P003_XACCXOR/Xdffa0/M9_d
+ N_XACCXOR/XDFFA0/N1_XACCXOR/Xdffa0/M9_g N_GND_XACCXOR/Xdffa0/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXACCXOR/Xdffa3/M9 N_XACCXOR/XDFFA3/P003_XACCXOR/Xdffa3/M9_d
+ N_XACCXOR/XDFFA3/N1_XACCXOR/Xdffa3/M9_g N_GND_XACCXOR/Xdffa3/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXACCXOR/Xdffa5/M9 N_XACCXOR/XDFFA5/P003_XACCXOR/Xdffa5/M9_d
+ N_XACCXOR/XDFFA5/N1_XACCXOR/Xdffa5/M9_g N_GND_XACCXOR/Xdffa5/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXACCXOR/Xdffa7/M9 N_XACCXOR/XDFFA7/P003_XACCXOR/Xdffa7/M9_d
+ N_XACCXOR/XDFFA7/N1_XACCXOR/Xdffa7/M9_g N_GND_XACCXOR/Xdffa7/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXACCXOR/Xdffa9/M9 N_XACCXOR/XDFFA9/P003_XACCXOR/Xdffa9/M9_d
+ N_XACCXOR/XDFFA9/N1_XACCXOR/Xdffa9/M9_g N_GND_XACCXOR/Xdffa9/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXACCXOR/Xdffa11/M9 N_XACCXOR/XDFFA11/P003_XACCXOR/Xdffa11/M9_d
+ N_XACCXOR/XDFFA11/N1_XACCXOR/Xdffa11/M9_g N_GND_XACCXOR/Xdffa11/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXADDER/Xa11/Xyb3/M38 N_XADDER/XA11/XYB3/N008_XADDER/Xa11/Xyb3/M38_d
+ N_XADDER/G1_XADDER/Xa11/Xyb3/M38_g N_GND_XADDER/Xa11/Xyb3/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe2/M21 N_XBOOTH/XE2/N004_XBOOTH/Xe2/M21_d
+ N_XBOOTH/A_D[4]_XBOOTH/Xe2/M21_g N_A_D[3]_XBOOTH/Xe2/M21_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xe1/M21 N_XBOOTH/XE1/N004_XBOOTH/Xe1/M21_d
+ N_XBOOTH/A_D[2]_XBOOTH/Xe1/M21_g N_A_D[1]_XBOOTH/Xe1/M21_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xe0/M21 N_XBOOTH/XE0/N004_XBOOTH/Xe0/M21_d
+ N_XBOOTH/A_D[0]_XBOOTH/Xe0/M21_g N_GND_XBOOTH/Xe0/M21_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa62/Xao1/M10 N_XADDER/XA62/XAO1/N004_XADDER/Xa62/Xao1/M10_d
+ N_XADDER/P2_XADDER/Xa62/Xao1/M10_g N_GND_XADDER/Xa62/Xao1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.86e-13
+ PD=2.8e-07 PS=1.74e-06
mX02/xd23/M3 N_X02/XD23/N0_X02/xd23/M3_d N_OUT1[2]_X02/xd23/M3_g
+ N_GND_X02/xd23/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa0/M11 N_XACCXOR/DACC[0]_XACCXOR/Xdffa0/M11_d
+ N_XACCXOR/XDFFA0/N3_XACCXOR/Xdffa0/M11_g N_GND_XACCXOR/Xdffa0/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXACCXOR/Xdffa3/M11 N_XACCXOR/DACC[3]_XACCXOR/Xdffa3/M11_d
+ N_XACCXOR/XDFFA3/N3_XACCXOR/Xdffa3/M11_g N_GND_XACCXOR/Xdffa3/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXACCXOR/Xdffa5/M11 N_XACCXOR/DACC[5]_XACCXOR/Xdffa5/M11_d
+ N_XACCXOR/XDFFA5/N3_XACCXOR/Xdffa5/M11_g N_GND_XACCXOR/Xdffa5/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXACCXOR/Xdffa7/M11 N_XACCXOR/DACC[7]_XACCXOR/Xdffa7/M11_d
+ N_XACCXOR/XDFFA7/N3_XACCXOR/Xdffa7/M11_g N_GND_XACCXOR/Xdffa7/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXACCXOR/Xdffa9/M11 N_XACCXOR/DACC[9]_XACCXOR/Xdffa9/M11_d
+ N_XACCXOR/XDFFA9/N3_XACCXOR/Xdffa9/M11_g N_GND_XACCXOR/Xdffa9/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXACCXOR/Xdffa11/M11 N_XACCXOR/DACC[11]_XACCXOR/Xdffa11/M11_d
+ N_XACCXOR/XDFFA11/N3_XACCXOR/Xdffa11/M11_g N_GND_XACCXOR/Xdffa11/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXADDER/Xa62/Xao1/M9 N_XADDER/XA62/XAO1/N003_XADDER/Xa62/Xao1/M9_d
+ N_XADDER/GG1_XADDER/Xa62/Xao1/M9_g
+ N_XADDER/XA62/XAO1/N004_XADDER/Xa62/Xao1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14 PD=1.44e-06 PS=2.8e-07
mXADDER/Xa03/Xrb2/M1 N_XADDER/XA03/XRB2/N002_XADDER/Xa03/Xrb2/M1_d
+ N_C[2]_XADDER/Xa03/Xrb2/M1_g N_S[2]_XADDER/Xa03/Xrb2/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/Xdffmod/M3 N_XCSA/XDFFMOD/N0_XCSA/Xdffmod/M3_d N_DMODE_XCSA/Xdffmod/M3_g
+ N_GND_XCSA/Xdffmod/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa12/M3 N_XCSA/XDFFA12/N0_XCSA/Xdffa12/M3_d
+ N_XCSA/LV3_S[0]_XCSA/Xdffa12/M3_g N_GND_XCSA/Xdffa12/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd23/M6 N_X02/XD23/P002_X02/xd23/M6_d N_CLK_X02/xd23/M6_g
+ N_GND_X02/xd23/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXADDER/Xa11/Xyb3/Xor1/M16 N_XADDER/GG1_XADDER/Xa11/Xyb3/Xor1/M16_d
+ N_XADDER/XA11/XYB3/N008_XADDER/Xa11/Xyb3/Xor1/M16_g
+ N_GND_XADDER/Xa11/Xyb3/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xe2/M23 N_XBOOTH/S2_XBOOTH/Xe2/M23_d N_XBOOTH/XE2/N004_XBOOTH/Xe2/M23_g
+ N_GND_XBOOTH/Xe2/M23_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xe1/M23 N_XBOOTH/S1_XBOOTH/Xe1/M23_d N_XBOOTH/XE1/N004_XBOOTH/Xe1/M23_g
+ N_GND_XBOOTH/Xe1/M23_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xe0/M23 N_XBOOTH/S0_XBOOTH/Xe0/M23_d N_XBOOTH/XE0/N004_XBOOTH/Xe0/M23_g
+ N_GND_XBOOTH/Xe0/M23_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa03/Xrb2/M2 N_XADDER/XA03/XRB2/N002_XADDER/Xa03/Xrb2/M2_d
+ N_S[2]_XADDER/Xa03/Xrb2/M2_g N_C[2]_XADDER/Xa03/Xrb2/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mX02/xd23/M5 N_X02/XD23/N1_X02/xd23/M5_d N_X02/XD23/N0_X02/xd23/M5_g
+ N_X02/XD23/P002_X02/xd23/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffmod/M6 N_XCSA/XDFFMOD/P002_XCSA/Xdffmod/M6_d N_CLK_XCSA/Xdffmod/M6_g
+ N_GND_XCSA/Xdffmod/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/Xdffa12/M6 N_XCSA/XDFFA12/P002_XCSA/Xdffa12/M6_d N_CLK_XCSA/Xdffa12/M6_g
+ N_GND_XCSA/Xdffa12/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXADDER/Xa23/Xao1/M9 N_XADDER/XA23/XAO1/N003_XADDER/Xa23/Xao1/M9_d
+ N_XADDER/GG1_XADDER/Xa23/Xao1/M9_g
+ N_XADDER/XA23/XAO1/N004_XADDER/Xa23/Xao1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14 PD=1.44e-06 PS=2.8e-07
mXACCXOR/X_xor0/M2 N_XACCXOR/X_XOR0/N002_XACCXOR/X_xor0/M2_d
+ N_DMODE_XACCXOR/X_xor0/M2_g N_XACCXOR/DACC[0]_XACCXOR/X_xor0/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXACCXOR/X_xor3/M2 N_XACCXOR/X_XOR3/N002_XACCXOR/X_xor3/M2_d
+ N_DMODE_XACCXOR/X_xor3/M2_g N_XACCXOR/DACC[3]_XACCXOR/X_xor3/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXACCXOR/X_xor5/M2 N_XACCXOR/X_XOR5/N002_XACCXOR/X_xor5/M2_d
+ N_DMODE_XACCXOR/X_xor5/M2_g N_XACCXOR/DACC[5]_XACCXOR/X_xor5/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXACCXOR/X_xor7/M2 N_XACCXOR/X_XOR7/N002_XACCXOR/X_xor7/M2_d
+ N_DMODE_XACCXOR/X_xor7/M2_g N_XACCXOR/DACC[7]_XACCXOR/X_xor7/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXACCXOR/X_xor9/M2 N_XACCXOR/X_XOR9/N002_XACCXOR/X_xor9/M2_d
+ N_DMODE_XACCXOR/X_xor9/M2_g N_XACCXOR/DACC[9]_XACCXOR/X_xor9/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXACCXOR/X_xor11/M2 N_XACCXOR/X_XOR11/N002_XACCXOR/X_xor11/M2_d
+ N_DMODE_XACCXOR/X_xor11/M2_g N_XACCXOR/DACC[11]_XACCXOR/X_xor11/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/Xdffmod/M5 N_XCSA/XDFFMOD/N1_XCSA/Xdffmod/M5_d
+ N_XCSA/XDFFMOD/N0_XCSA/Xdffmod/M5_g N_XCSA/XDFFMOD/P002_XCSA/Xdffmod/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa12/M5 N_XCSA/XDFFA12/N1_XCSA/Xdffa12/M5_d
+ N_XCSA/XDFFA12/N0_XCSA/Xdffa12/M5_g N_XCSA/XDFFA12/P002_XCSA/Xdffa12/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa23/Xao1/M10 N_XADDER/XA23/XAO1/N004_XADDER/Xa23/Xao1/M10_d
+ N_XADDER/PP3_XADDER/Xa23/Xao1/M10_g N_GND_XADDER/Xa23/Xao1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.86e-13
+ PD=2.8e-07 PS=1.74e-06
mXACCXOR/X_xor0/M1 N_XACCXOR/X_XOR0/N002_XACCXOR/X_xor0/M1_d
+ N_XACCXOR/DACC[0]_XACCXOR/X_xor0/M1_g N_DMODE_XACCXOR/X_xor0/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXACCXOR/X_xor3/M1 N_XACCXOR/X_XOR3/N002_XACCXOR/X_xor3/M1_d
+ N_XACCXOR/DACC[3]_XACCXOR/X_xor3/M1_g N_DMODE_XACCXOR/X_xor3/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXACCXOR/X_xor5/M1 N_XACCXOR/X_XOR5/N002_XACCXOR/X_xor5/M1_d
+ N_XACCXOR/DACC[5]_XACCXOR/X_xor5/M1_g N_DMODE_XACCXOR/X_xor5/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXACCXOR/X_xor7/M1 N_XACCXOR/X_XOR7/N002_XACCXOR/X_xor7/M1_d
+ N_XACCXOR/DACC[7]_XACCXOR/X_xor7/M1_g N_DMODE_XACCXOR/X_xor7/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXACCXOR/X_xor9/M1 N_XACCXOR/X_XOR9/N002_XACCXOR/X_xor9/M1_d
+ N_XACCXOR/DACC[9]_XACCXOR/X_xor9/M1_g N_DMODE_XACCXOR/X_xor9/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXACCXOR/X_xor11/M1 N_XACCXOR/X_XOR11/N002_XACCXOR/X_xor11/M1_d
+ N_XACCXOR/DACC[11]_XACCXOR/X_xor11/M1_g N_DMODE_XACCXOR/X_xor11/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa13/Xyb1/Xand1/M16 N_XADDER/PP3_XADDER/Xa13/Xyb1/Xand1/M16_d
+ N_XADDER/XA13/XYB1/N003_XADDER/Xa13/Xyb1/Xand1/M16_g
+ N_GND_XADDER/Xa13/Xyb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd23/M8 N_X02/XD23/N3_X02/xd23/M8_d N_CLK_X02/xd23/M8_g
+ N_X02/XD23/P003_X02/xd23/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa03/Xrb1/M10 N_XADDER/XA03/XRB1/N004_XADDER/Xa03/Xrb1/M10_d
+ N_S[2]_XADDER/Xa03/Xrb1/M10_g N_GND_XADDER/Xa03/Xrb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXBOOTH/Xsel20/M2 N_noxref_2105_XBOOTH/Xsel20/M2_d N_GND_XBOOTH/Xsel20/M2_g
+ N_GND_XBOOTH/Xsel20/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel10/M2 N_noxref_2106_XBOOTH/Xsel10/M2_d N_GND_XBOOTH/Xsel10/M2_g
+ N_GND_XBOOTH/Xsel10/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel00/M2 N_noxref_2107_XBOOTH/Xsel00/M2_d N_GND_XBOOTH/Xsel00/M2_g
+ N_GND_XBOOTH/Xsel00/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mX02/xd23/M9 N_X02/XD23/P003_X02/xd23/M9_d N_X02/XD23/N1_X02/xd23/M9_g
+ N_GND_X02/xd23/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.76e-13 PD=2.8e-07 PS=8e-07
mXADDER/Xa03/Xrb1/M9 N_XADDER/XA03/XRB1/N003_XADDER/Xa03/Xrb1/M9_d
+ N_C[2]_XADDER/Xa03/Xrb1/M9_g N_XADDER/XA03/XRB1/N004_XADDER/Xa03/Xrb1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14
+ PD=1.44e-06 PS=2.8e-07
mXCSA/Xdffmod/M8 N_XCSA/XDFFMOD/N3_XCSA/Xdffmod/M8_d N_CLK_XCSA/Xdffmod/M8_g
+ N_XCSA/XDFFMOD/P003_XCSA/Xdffmod/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa12/M8 N_XCSA/XDFFA12/N3_XCSA/Xdffa12/M8_d N_CLK_XCSA/Xdffa12/M8_g
+ N_XCSA/XDFFA12/P003_XCSA/Xdffa12/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel20/M1 N_XBOOTH/XSEL20/N002_XBOOTH/Xsel20/M1_d
+ N_XBOOTH/D2_XBOOTH/Xsel20/M1_g N_noxref_2105_XBOOTH/Xsel20/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel10/M1 N_XBOOTH/XSEL10/N002_XBOOTH/Xsel10/M1_d
+ N_XBOOTH/D1_XBOOTH/Xsel10/M1_g N_noxref_2106_XBOOTH/Xsel10/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel00/M1 N_XBOOTH/XSEL00/N002_XBOOTH/Xsel00/M1_d
+ N_XBOOTH/D0_XBOOTH/Xsel00/M1_g N_noxref_2107_XBOOTH/Xsel00/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXCSA/Xdffmod/M9 N_XCSA/XDFFMOD/P003_XCSA/Xdffmod/M9_d
+ N_XCSA/XDFFMOD/N1_XCSA/Xdffmod/M9_g N_GND_XCSA/Xdffmod/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXADDER/Xa23/Xao1/Xand1/M16 N_XADDER/XA23/OUT1_XADDER/Xa23/Xao1/Xand1/M16_d
+ N_XADDER/XA23/XAO1/N003_XADDER/Xa23/Xao1/Xand1/M16_g
+ N_GND_XADDER/Xa23/Xao1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa12/M9 N_XCSA/XDFFA12/P003_XCSA/Xdffa12/M9_d
+ N_XCSA/XDFFA12/N1_XCSA/Xdffa12/M9_g N_GND_XCSA/Xdffa12/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXACCXOR/X_xor0/M3 N_CACC[0]_XACCXOR/X_xor0/M3_d
+ N_XACCXOR/X_XOR0/N002_XACCXOR/X_xor0/M3_g N_GND_XACCXOR/X_xor0/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor3/M3 N_CACC[3]_XACCXOR/X_xor3/M3_d
+ N_XACCXOR/X_XOR3/N002_XACCXOR/X_xor3/M3_g N_GND_XACCXOR/X_xor3/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor5/M3 N_CACC[5]_XACCXOR/X_xor5/M3_d
+ N_XACCXOR/X_XOR5/N002_XACCXOR/X_xor5/M3_g N_GND_XACCXOR/X_xor5/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor7/M3 N_CACC[7]_XACCXOR/X_xor7/M3_d
+ N_XACCXOR/X_XOR7/N002_XACCXOR/X_xor7/M3_g N_GND_XACCXOR/X_xor7/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor9/M3 N_CACC[9]_XACCXOR/X_xor9/M3_d
+ N_XACCXOR/X_XOR9/N002_XACCXOR/X_xor9/M3_g N_GND_XACCXOR/X_xor9/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor11/M3 N_CACC[11]_XACCXOR/X_xor11/M3_d
+ N_XACCXOR/X_XOR11/N002_XACCXOR/X_xor11/M3_g N_GND_XACCXOR/X_xor11/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa13/Xyb1/M9 N_XADDER/XA13/XYB1/N003_XADDER/Xa13/Xyb1/M9_d
+ N_XADDER/P2_XADDER/Xa13/Xyb1/M9_g
+ N_XADDER/XA13/XYB1/N004_XADDER/Xa13/Xyb1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=9.24e-14 PD=1.44e-06 PS=4.2e-07
mX02/xd23/M11 N_OUT[2]_X02/xd23/M11_d N_X02/XD23/N3_X02/xd23/M11_g
+ N_GND_X02/xd23/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXBOOTH/Xsel20/M3 N_XBOOTH/XSEL20/N002_XBOOTH/Xsel20/M3_d
+ N_XBOOTH/S2_XBOOTH/Xsel20/M3_g N_noxref_2111_XBOOTH/Xsel20/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel10/M3 N_XBOOTH/XSEL10/N002_XBOOTH/Xsel10/M3_d
+ N_XBOOTH/S1_XBOOTH/Xsel10/M3_g N_noxref_2112_XBOOTH/Xsel10/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel00/M3 N_XBOOTH/XSEL00/N002_XBOOTH/Xsel00/M3_d
+ N_XBOOTH/S0_XBOOTH/Xsel00/M3_g N_noxref_2113_XBOOTH/Xsel00/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXADDER/Xa13/Xyb1/M10 N_XADDER/XA13/XYB1/N004_XADDER/Xa13/Xyb1/M10_d
+ N_XADDER/P3_XADDER/Xa13/Xyb1/M10_g N_GND_XADDER/Xa13/Xyb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=9.24e-14 AS=2.244e-13
+ PD=4.2e-07 PS=1.46e-06
mXADDER/Xa03/Xrb1/Xand1/M16 N_XADDER/G2_XADDER/Xa03/Xrb1/Xand1/M16_d
+ N_XADDER/XA03/XRB1/N003_XADDER/Xa03/Xrb1/Xand1/M16_g
+ N_GND_XADDER/Xa03/Xrb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffmod/M11 N_CIN_XCSA/Xdffmod/M11_d N_XCSA/XDFFMOD/N3_XCSA/Xdffmod/M11_g
+ N_GND_XCSA/Xdffmod/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/Xdffa12/M11 N_S[0]_XCSA/Xdffa12/M11_d N_XCSA/XDFFA12/N3_XCSA/Xdffa12/M11_g
+ N_GND_XCSA/Xdffa12/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXBOOTH/Xsel20/M4 N_noxref_2111_XBOOTH/Xsel20/M4_d
+ N_XBOOTH/B_D[0]_XBOOTH/Xsel20/M4_g N_GND_XBOOTH/Xsel20/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel10/M4 N_noxref_2112_XBOOTH/Xsel10/M4_d
+ N_XBOOTH/B_D[0]_XBOOTH/Xsel10/M4_g N_GND_XBOOTH/Xsel10/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel00/M4 N_noxref_2113_XBOOTH/Xsel00/M4_d
+ N_XBOOTH/B_D[0]_XBOOTH/Xsel00/M4_g N_GND_XBOOTH/Xsel00/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXADDER/Xa23/Xao2/M37 N_XADDER/XA23/XAO2/N008_XADDER/Xa23/Xao2/M37_d
+ N_XADDER/XA23/OUT1_XADDER/Xa23/Xao2/M37_g N_GND_XADDER/Xa23/Xao2/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xdffb0/M3 N_XBOOTH/XDFFB0/N0_XBOOTH/Xdffb0/M3_d
+ N_B[0]_XBOOTH/Xdffb0/M3_g N_GND_XBOOTH/Xdffb0/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd24/M3 N_X02/XD24/N0_X02/xd24/M3_d N_OUT1[3]_X02/xd24/M3_g
+ N_GND_X02/xd24/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_HA0/M14 N_XCSA/LV1_C[3]_XCSA/X_LV1_HA0/M14_d
+ N_XCSA/X_LV1_HA0/N001_XCSA/X_LV1_HA0/M14_g N_GND_XCSA/X_LV1_HA0/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_HA0/X_xor/M3 N_XCSA/LV1_S[2]_XCSA/X_LV1_HA0/X_xor/M3_d
+ N_XCSA/X_LV1_HA0/X_XOR/N002_XCSA/X_LV1_HA0/X_xor/M3_g
+ N_GND_XCSA/X_LV1_HA0/X_xor/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel20/M5 N_XBOOTH/XSEL20/B_XBOOTH/Xsel20/M5_d
+ N_XBOOTH/XSEL20/N002_XBOOTH/Xsel20/M5_g N_GND_XBOOTH/Xsel20/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel10/M5 N_XBOOTH/XSEL10/B_XBOOTH/Xsel10/M5_d
+ N_XBOOTH/XSEL10/N002_XBOOTH/Xsel10/M5_g N_GND_XBOOTH/Xsel10/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel00/M5 N_XBOOTH/XSEL00/B_XBOOTH/Xsel00/M5_d
+ N_XBOOTH/XSEL00/N002_XBOOTH/Xsel00/M5_g N_GND_XBOOTH/Xsel00/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa23/Xao2/M38 N_XADDER/XA23/XAO2/N008_XADDER/Xa23/Xao2/M38_d
+ N_XADDER/GG3_XADDER/Xa23/Xao2/M38_g N_GND_XADDER/Xa23/Xao2/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xdffb0/M6 N_XBOOTH/XDFFB0/P002_XBOOTH/Xdffb0/M6_d
+ N_CLK_XBOOTH/Xdffb0/M6_g N_GND_XBOOTH/Xdffb0/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXADDER/Xa13/Xyb2/M10 N_XADDER/XA13/XYB2/N004_XADDER/Xa13/Xyb2/M10_d
+ N_XADDER/P3_XADDER/Xa13/Xyb2/M10_g N_GND_XADDER/Xa13/Xyb2/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXCSA/Xdffa0/M3 N_XCSA/XDFFA0/N0_XCSA/Xdffa0/M3_d
+ N_XCSA/LV3_C[1]_XCSA/Xdffa0/M3_g N_GND_XCSA/Xdffa0/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa13/M3 N_XCSA/XDFFA13/N0_XCSA/Xdffa13/M3_d
+ N_XCSA/LV3_S[1]_XCSA/Xdffa13/M3_g N_GND_XCSA/Xdffa13/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd24/M6 N_X02/XD24/P002_X02/xd24/M6_d N_CLK_X02/xd24/M6_g
+ N_GND_X02/xd24/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/X_LV2_HA1/X_xor/M1 N_XCSA/X_LV2_HA1/X_XOR/N002_XCSA/X_LV2_HA1/X_xor/M1_d
+ N_A_D[3]_XCSA/X_LV2_HA1/X_xor/M1_g N_XCSA/LV1_S[2]_XCSA/X_LV2_HA1/X_xor/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA1/M12 N_XCSA/X_LV2_HA1/P001_XCSA/X_LV2_HA1/M12_d
+ N_A_D[3]_XCSA/X_LV2_HA1/M12_g N_GND_XCSA/X_LV2_HA1/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXADDER/Xa04/Xrb2/M3 N_XADDER/P3_XADDER/Xa04/Xrb2/M3_d
+ N_XADDER/XA04/XRB2/N002_XADDER/Xa04/Xrb2/M3_g N_GND_XADDER/Xa04/Xrb2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xdffb0/M5 N_XBOOTH/XDFFB0/N1_XBOOTH/Xdffb0/M5_d
+ N_XBOOTH/XDFFB0/N0_XBOOTH/Xdffb0/M5_g N_XBOOTH/XDFFB0/P002_XBOOTH/Xdffb0/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa13/Xyb2/M9 N_XADDER/XA13/XYB2/N003_XADDER/Xa13/Xyb2/M9_d
+ N_XADDER/G2_XADDER/Xa13/Xyb2/M9_g
+ N_XADDER/XA13/XYB2/N004_XADDER/Xa13/Xyb2/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=6.16e-14 PD=1.74e-06 PS=2.8e-07
mX02/xd24/M5 N_X02/XD24/N1_X02/xd24/M5_d N_X02/XD24/N0_X02/xd24/M5_g
+ N_X02/XD24/P002_X02/xd24/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV3_HA0/M11 N_XCSA/X_LV3_HA0/P001_XCSA/X_LV3_HA0/M11_d
+ N_XCSA/LV2_S[0]_XCSA/X_LV3_HA0/M11_g N_GND_XCSA/X_LV3_HA0/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV3_HA0/X_xor/M2 N_XCSA/X_LV3_HA0/X_XOR/N002_XCSA/X_LV3_HA0/X_xor/M2_d
+ N_XCSA/LV2_S[0]_XCSA/X_LV3_HA0/X_xor/M2_g N_CACC[0]_XCSA/X_LV3_HA0/X_xor/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/Xdffa0/M6 N_XCSA/XDFFA0/P002_XCSA/Xdffa0/M6_d N_CLK_XCSA/Xdffa0/M6_g
+ N_GND_XCSA/Xdffa0/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/Xdffa13/M6 N_XCSA/XDFFA13/P002_XCSA/Xdffa13/M6_d N_CLK_XCSA/Xdffa13/M6_g
+ N_GND_XCSA/Xdffa13/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/X_LV2_HA1/X_xor/M2 N_XCSA/X_LV2_HA1/X_XOR/N002_XCSA/X_LV2_HA1/X_xor/M2_d
+ N_XCSA/LV1_S[2]_XCSA/X_LV2_HA1/X_xor/M2_g N_A_D[3]_XCSA/X_LV2_HA1/X_xor/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_HA1/M11 N_XCSA/X_LV2_HA1/N001_XCSA/X_LV2_HA1/M11_d
+ N_XCSA/LV1_S[2]_XCSA/X_LV2_HA1/M11_g
+ N_XCSA/X_LV2_HA1/P001_XCSA/X_LV2_HA1/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_HA0/M12 N_XCSA/X_LV1_HA0/N001_XCSA/X_LV1_HA0/M12_d
+ N_PP1[0]_XCSA/X_LV1_HA0/M12_g N_XCSA/X_LV1_HA0/P001_XCSA/X_LV1_HA0/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_HA0/X_xor/M1 N_XCSA/X_LV1_HA0/X_XOR/N002_XCSA/X_LV1_HA0/X_xor/M1_d
+ N_PP1[0]_XCSA/X_LV1_HA0/X_xor/M1_g N_PP0[2]_XCSA/X_LV1_HA0/X_xor/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/Xdffa0/M5 N_XCSA/XDFFA0/N1_XCSA/Xdffa0/M5_d
+ N_XCSA/XDFFA0/N0_XCSA/Xdffa0/M5_g N_XCSA/XDFFA0/P002_XCSA/Xdffa0/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa23/Xao2/Xor1/M16 N_XADDER/GGG3_XADDER/Xa23/Xao2/Xor1/M16_d
+ N_XADDER/XA23/XAO2/N008_XADDER/Xa23/Xao2/Xor1/M16_g
+ N_GND_XADDER/Xa23/Xao2/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa13/M5 N_XCSA/XDFFA13/N1_XCSA/Xdffa13/M5_d
+ N_XCSA/XDFFA13/N0_XCSA/Xdffa13/M5_g N_XCSA/XDFFA13/P002_XCSA/Xdffa13/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV3_HA0/M12 N_XCSA/X_LV3_HA0/N001_XCSA/X_LV3_HA0/M12_d
+ N_CACC[0]_XCSA/X_LV3_HA0/M12_g N_XCSA/X_LV3_HA0/P001_XCSA/X_LV3_HA0/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_HA0/X_xor/M1 N_XCSA/X_LV3_HA0/X_XOR/N002_XCSA/X_LV3_HA0/X_xor/M1_d
+ N_CACC[0]_XCSA/X_LV3_HA0/X_xor/M1_g N_XCSA/LV2_S[0]_XCSA/X_LV3_HA0/X_xor/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa04/Xrb2/M1 N_XADDER/XA04/XRB2/N002_XADDER/Xa04/Xrb2/M1_d
+ N_C[3]_XADDER/Xa04/Xrb2/M1_g N_S[3]_XADDER/Xa04/Xrb2/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel20/M12 N_XBOOTH/XSEL20/N004_XBOOTH/Xsel20/M12_d
+ N_A_D[5]_XBOOTH/Xsel20/M12_g N_XBOOTH/XSEL20/B_XBOOTH/Xsel20/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel10/M12 N_XBOOTH/XSEL10/N004_XBOOTH/Xsel10/M12_d
+ N_A_D[3]_XBOOTH/Xsel10/M12_g N_XBOOTH/XSEL10/B_XBOOTH/Xsel10/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel00/M12 N_XBOOTH/XSEL00/N004_XBOOTH/Xsel00/M12_d
+ N_A_D[1]_XBOOTH/Xsel00/M12_g N_XBOOTH/XSEL00/B_XBOOTH/Xsel00/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xdffb0/M8 N_XBOOTH/XDFFB0/N3_XBOOTH/Xdffb0/M8_d N_CLK_XBOOTH/Xdffb0/M8_g
+ N_XBOOTH/XDFFB0/P003_XBOOTH/Xdffb0/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV1_HA0/M11 N_XCSA/X_LV1_HA0/P001_XCSA/X_LV1_HA0/M11_d
+ N_PP0[2]_XCSA/X_LV1_HA0/M11_g N_GND_XCSA/X_LV1_HA0/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV1_HA0/X_xor/M2 N_XCSA/X_LV1_HA0/X_XOR/N002_XCSA/X_LV1_HA0/X_xor/M2_d
+ N_PP0[2]_XCSA/X_LV1_HA0/X_xor/M2_g N_PP1[0]_XCSA/X_LV1_HA0/X_xor/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXADDER/Xa13/Xyb2/Xand1/M16 N_XADDER/XA13/T1_XADDER/Xa13/Xyb2/Xand1/M16_d
+ N_XADDER/XA13/XYB2/N003_XADDER/Xa13/Xyb2/Xand1/M16_g
+ N_GND_XADDER/Xa13/Xyb2/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd24/M8 N_X02/XD24/N3_X02/xd24/M8_d N_CLK_X02/xd24/M8_g
+ N_X02/XD24/P003_X02/xd24/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xdffb0/M9 N_XBOOTH/XDFFB0/P003_XBOOTH/Xdffb0/M9_d
+ N_XBOOTH/XDFFB0/N1_XBOOTH/Xdffb0/M9_g N_GND_XBOOTH/Xdffb0/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/X_LV2_HA1/X_xor/M3 N_XCSA/LV2_S[2]_XCSA/X_LV2_HA1/X_xor/M3_d
+ N_XCSA/X_LV2_HA1/X_XOR/N002_XCSA/X_LV2_HA1/X_xor/M3_g
+ N_GND_XCSA/X_LV2_HA1/X_xor/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA1/M14 N_XCSA/LV2_C[3]_XCSA/X_LV2_HA1/M14_d
+ N_XCSA/X_LV2_HA1/N001_XCSA/X_LV2_HA1/M14_g N_GND_XCSA/X_LV2_HA1/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa04/Xrb2/M2 N_XADDER/XA04/XRB2/N002_XADDER/Xa04/Xrb2/M2_d
+ N_S[3]_XADDER/Xa04/Xrb2/M2_g N_C[3]_XADDER/Xa04/Xrb2/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mX02/xd24/M9 N_X02/XD24/P003_X02/xd24/M9_d N_X02/XD24/N1_X02/xd24/M9_g
+ N_GND_X02/xd24/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.76e-13 PD=2.8e-07 PS=8e-07
mXBOOTH/Xsel20/M11 N_XBOOTH/XSEL20/N004_XBOOTH/Xsel20/M11_d
+ N_XBOOTH/XSEL20/B_XBOOTH/Xsel20/M11_g N_A_D[5]_XBOOTH/Xsel20/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel10/M11 N_XBOOTH/XSEL10/N004_XBOOTH/Xsel10/M11_d
+ N_XBOOTH/XSEL10/B_XBOOTH/Xsel10/M11_g N_A_D[3]_XBOOTH/Xsel10/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel00/M11 N_XBOOTH/XSEL00/N004_XBOOTH/Xsel00/M11_d
+ N_XBOOTH/XSEL00/B_XBOOTH/Xsel00/M11_g N_A_D[1]_XBOOTH/Xsel00/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/Xdffa0/M8 N_XCSA/XDFFA0/N3_XCSA/Xdffa0/M8_d N_CLK_XCSA/Xdffa0/M8_g
+ N_XCSA/XDFFA0/P003_XCSA/Xdffa0/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa13/M8 N_XCSA/XDFFA13/N3_XCSA/Xdffa13/M8_d N_CLK_XCSA/Xdffa13/M8_g
+ N_XCSA/XDFFA13/P003_XCSA/Xdffa13/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa55/Xao1/M9 N_XADDER/XA55/XAO1/N003_XADDER/Xa55/Xao1/M9_d
+ N_XADDER/GGG3_XADDER/Xa55/Xao1/M9_g
+ N_XADDER/XA55/XAO1/N004_XADDER/Xa55/Xao1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14 PD=1.44e-06 PS=2.8e-07
mXCSA/X_LV3_HA0/M14 N_XCSA/LV3_C[1]_XCSA/X_LV3_HA0/M14_d
+ N_XCSA/X_LV3_HA0/N001_XCSA/X_LV3_HA0/M14_g N_GND_XCSA/X_LV3_HA0/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_HA0/X_xor/M3 N_XCSA/LV3_S[0]_XCSA/X_LV3_HA0/X_xor/M3_d
+ N_XCSA/X_LV3_HA0/X_XOR/N002_XCSA/X_LV3_HA0/X_xor/M3_g
+ N_GND_XCSA/X_LV3_HA0/X_xor/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa0/M9 N_XCSA/XDFFA0/P003_XCSA/Xdffa0/M9_d
+ N_XCSA/XDFFA0/N1_XCSA/Xdffa0/M9_g N_GND_XCSA/Xdffa0/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/Xdffa13/M9 N_XCSA/XDFFA13/P003_XCSA/Xdffa13/M9_d
+ N_XCSA/XDFFA13/N1_XCSA/Xdffa13/M9_g N_GND_XCSA/Xdffa13/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXADDER/Xa55/Xao1/M10 N_XADDER/XA55/XAO1/N004_XADDER/Xa55/Xao1/M10_d
+ N_XADDER/PP5_XADDER/Xa55/Xao1/M10_g N_GND_XADDER/Xa55/Xao1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.86e-13
+ PD=2.8e-07 PS=1.74e-06
mXBOOTH/Xdffb0/M11 N_XBOOTH/B_D[0]_XBOOTH/Xdffb0/M11_d
+ N_XBOOTH/XDFFB0/N3_XBOOTH/Xdffb0/M11_g N_GND_XBOOTH/Xdffb0/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXADDER/Xa13/Xyb3/M37 N_XADDER/XA13/XYB3/N008_XADDER/Xa13/Xyb3/M37_d
+ N_XADDER/XA13/T1_XADDER/Xa13/Xyb3/M37_g N_GND_XADDER/Xa13/Xyb3/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd24/M11 N_OUT[3]_X02/xd24/M11_d N_X02/XD24/N3_X02/xd24/M11_g
+ N_GND_X02/xd24/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXBOOTH/Xsel20/M13 N_PP2[0]_XBOOTH/Xsel20/M13_d
+ N_XBOOTH/XSEL20/N004_XBOOTH/Xsel20/M13_g N_GND_XBOOTH/Xsel20/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel10/M13 N_PP1[0]_XBOOTH/Xsel10/M13_d
+ N_XBOOTH/XSEL10/N004_XBOOTH/Xsel10/M13_g N_GND_XBOOTH/Xsel10/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel00/M13 N_PP0[0]_XBOOTH/Xsel00/M13_d
+ N_XBOOTH/XSEL00/N004_XBOOTH/Xsel00/M13_g N_GND_XBOOTH/Xsel00/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa04/Xrb1/M10 N_XADDER/XA04/XRB1/N004_XADDER/Xa04/Xrb1/M10_d
+ N_S[3]_XADDER/Xa04/Xrb1/M10_g N_GND_XADDER/Xa04/Xrb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXCSA/Xdffa0/M11 N_C[1]_XCSA/Xdffa0/M11_d N_XCSA/XDFFA0/N3_XCSA/Xdffa0/M11_g
+ N_GND_XCSA/Xdffa0/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/Xdffa13/M11 N_S[1]_XCSA/Xdffa13/M11_d N_XCSA/XDFFA13/N3_XCSA/Xdffa13/M11_g
+ N_GND_XCSA/Xdffa13/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXADDER/Xa13/Xyb3/M38 N_XADDER/XA13/XYB3/N008_XADDER/Xa13/Xyb3/M38_d
+ N_XADDER/G3_XADDER/Xa13/Xyb3/M38_g N_GND_XADDER/Xa13/Xyb3/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_HA1/M14 N_XCSA/LV1_C[4]_XCSA/X_LV1_HA1/M14_d
+ N_XCSA/X_LV1_HA1/N001_XCSA/X_LV1_HA1/M14_g N_GND_XCSA/X_LV1_HA1/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_HA1/X_xor/M3 N_XCSA/LV1_S[3]_XCSA/X_LV1_HA1/X_xor/M3_d
+ N_XCSA/X_LV1_HA1/X_XOR/N002_XCSA/X_LV1_HA1/X_xor/M3_g
+ N_GND_XCSA/X_LV1_HA1/X_xor/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa04/Xrb1/M9 N_XADDER/XA04/XRB1/N003_XADDER/Xa04/Xrb1/M9_d
+ N_C[3]_XADDER/Xa04/Xrb1/M9_g N_XADDER/XA04/XRB1/N004_XADDER/Xa04/Xrb1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14
+ PD=1.44e-06 PS=2.8e-07
mXCSA/X_LV2_HA2/X_xor/M2 N_XCSA/X_LV2_HA2/X_XOR/N002_XCSA/X_LV2_HA2/X_xor/M2_d
+ N_XCSA/LV1_C[3]_XCSA/X_LV2_HA2/X_xor/M2_g
+ N_XCSA/LV1_S[3]_XCSA/X_LV2_HA2/X_xor/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13 PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA2/M11 N_XCSA/X_LV2_HA2/P001_XCSA/X_LV2_HA2/M11_d
+ N_XCSA/LV1_C[3]_XCSA/X_LV2_HA2/M11_g N_GND_XCSA/X_LV2_HA2/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXADDER/Xa55/Xao1/Xand1/M16 N_XADDER/XA55/OUT1_XADDER/Xa55/Xao1/Xand1/M16_d
+ N_XADDER/XA55/XAO1/N003_XADDER/Xa55/Xao1/Xand1/M16_g
+ N_GND_XADDER/Xa55/Xao1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA0/M25 N_XCSA/LV3_S[1]_XCSA/X_LV3_FA0/M25_d
+ N_XCSA/X_LV3_FA0/_SUM_XCSA/X_LV3_FA0/M25_g N_GND_XCSA/X_LV3_FA0/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.244e-13 AS=2.156e-13
+ PD=1.46e-06 PS=1.42e-06
mX02/xd25/M3 N_X02/XD25/N0_X02/xd25/M3_d N_OUT1[4]_X02/xd25/M3_g
+ N_GND_X02/xd25/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV2_HA2/X_xor/M1 N_XCSA/X_LV2_HA2/X_XOR/N002_XCSA/X_LV2_HA2/X_xor/M1_d
+ N_XCSA/LV1_S[3]_XCSA/X_LV2_HA2/X_xor/M1_g
+ N_XCSA/LV1_C[3]_XCSA/X_LV2_HA2/X_xor/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_HA2/M12 N_XCSA/X_LV2_HA2/N001_XCSA/X_LV2_HA2/M12_d
+ N_XCSA/LV1_S[3]_XCSA/X_LV2_HA2/M12_g
+ N_XCSA/X_LV2_HA2/P001_XCSA/X_LV2_HA2/M12_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa1/M3 N_XCSA/XDFFA1/N0_XCSA/Xdffa1/M3_d
+ N_XCSA/LV3_C[2]_XCSA/Xdffa1/M3_g N_GND_XCSA/Xdffa1/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa14/M3 N_XCSA/XDFFA14/N0_XCSA/Xdffa14/M3_d
+ N_XCSA/LV3_S[2]_XCSA/Xdffa14/M3_g N_GND_XCSA/Xdffa14/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa13/Xyb3/Xor1/M16 N_XADDER/GG3_XADDER/Xa13/Xyb3/Xor1/M16_d
+ N_XADDER/XA13/XYB3/N008_XADDER/Xa13/Xyb3/Xor1/M16_g
+ N_GND_XADDER/Xa13/Xyb3/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd25/M6 N_X02/XD25/P002_X02/xd25/M6_d N_CLK_X02/xd25/M6_g
+ N_GND_X02/xd25/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/X_LV3_FA0/M26 N_XCSA/LV3_C[2]_XCSA/X_LV3_FA0/M26_d
+ N_XCSA/X_LV3_FA0/_COUT_XCSA/X_LV3_FA0/M26_g N_GND_XCSA/X_LV3_FA0/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_HA1/M12 N_XCSA/X_LV1_HA1/N001_XCSA/X_LV1_HA1/M12_d
+ N_PP1[1]_XCSA/X_LV1_HA1/M12_g N_XCSA/X_LV1_HA1/P001_XCSA/X_LV1_HA1/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_HA1/X_xor/M1 N_XCSA/X_LV1_HA1/X_XOR/N002_XCSA/X_LV1_HA1/X_xor/M1_d
+ N_PP1[1]_XCSA/X_LV1_HA1/X_xor/M1_g N_PP0[3]_XCSA/X_LV1_HA1/X_xor/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel21/M2 N_noxref_2131_XBOOTH/Xsel21/M2_d
+ N_XBOOTH/B_D[0]_XBOOTH/Xsel21/M2_g N_GND_XBOOTH/Xsel21/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel11/M2 N_noxref_2132_XBOOTH/Xsel11/M2_d
+ N_XBOOTH/B_D[0]_XBOOTH/Xsel11/M2_g N_GND_XBOOTH/Xsel11/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel01/M2 N_noxref_2133_XBOOTH/Xsel01/M2_d
+ N_XBOOTH/B_D[0]_XBOOTH/Xsel01/M2_g N_GND_XBOOTH/Xsel01/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa04/Xrb1/Xand1/M16 N_XADDER/G3_XADDER/Xa04/Xrb1/Xand1/M16_d
+ N_XADDER/XA04/XRB1/N003_XADDER/Xa04/Xrb1/Xand1/M16_g
+ N_GND_XADDER/Xa04/Xrb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd25/M5 N_X02/XD25/N1_X02/xd25/M5_d N_X02/XD25/N0_X02/xd25/M5_g
+ N_X02/XD25/P002_X02/xd25/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa55/Xao2/M37 N_XADDER/XA55/XAO2/N008_XADDER/Xa55/Xao2/M37_d
+ N_XADDER/XA55/OUT1_XADDER/Xa55/Xao2/M37_g N_GND_XADDER/Xa55/Xao2/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA0/M21 N_XCSA/X_LV3_FA0/_SUM_XCSA/X_LV3_FA0/M21_d
+ N_XCSA/X_LV3_FA0/_COUT_XCSA/X_LV3_FA0/M21_g
+ N_XCSA/X_LV3_FA0/N004_XCSA/X_LV3_FA0/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXCSA/Xdffa1/M6 N_XCSA/XDFFA1/P002_XCSA/Xdffa1/M6_d N_CLK_XCSA/Xdffa1/M6_g
+ N_GND_XCSA/Xdffa1/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/Xdffa14/M6 N_XCSA/XDFFA14/P002_XCSA/Xdffa14/M6_d N_CLK_XCSA/Xdffa14/M6_g
+ N_GND_XCSA/Xdffa14/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/X_LV1_HA1/M11 N_XCSA/X_LV1_HA1/P001_XCSA/X_LV1_HA1/M11_d
+ N_PP0[3]_XCSA/X_LV1_HA1/M11_g N_GND_XCSA/X_LV1_HA1/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV1_HA1/X_xor/M2 N_XCSA/X_LV1_HA1/X_XOR/N002_XCSA/X_LV1_HA1/X_xor/M2_d
+ N_PP0[3]_XCSA/X_LV1_HA1/X_xor/M2_g N_PP1[1]_XCSA/X_LV1_HA1/X_xor/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXBOOTH/Xsel21/M1 N_XBOOTH/XSEL21/N002_XBOOTH/Xsel21/M1_d
+ N_XBOOTH/D2_XBOOTH/Xsel21/M1_g N_noxref_2131_XBOOTH/Xsel21/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel11/M1 N_XBOOTH/XSEL11/N002_XBOOTH/Xsel11/M1_d
+ N_XBOOTH/D1_XBOOTH/Xsel11/M1_g N_noxref_2132_XBOOTH/Xsel11/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel01/M1 N_XBOOTH/XSEL01/N002_XBOOTH/Xsel01/M1_d
+ N_XBOOTH/D0_XBOOTH/Xsel01/M1_g N_noxref_2133_XBOOTH/Xsel01/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXCSA/Xdffa1/M5 N_XCSA/XDFFA1/N1_XCSA/Xdffa1/M5_d
+ N_XCSA/XDFFA1/N0_XCSA/Xdffa1/M5_g N_XCSA/XDFFA1/P002_XCSA/Xdffa1/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa14/M5 N_XCSA/XDFFA14/N1_XCSA/Xdffa14/M5_d
+ N_XCSA/XDFFA14/N0_XCSA/Xdffa14/M5_g N_XCSA/XDFFA14/P002_XCSA/Xdffa14/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV2_HA2/X_xor/M3 N_XCSA/LV2_S[3]_XCSA/X_LV2_HA2/X_xor/M3_d
+ N_XCSA/X_LV2_HA2/X_XOR/N002_XCSA/X_LV2_HA2/X_xor/M3_g
+ N_GND_XCSA/X_LV2_HA2/X_xor/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA2/M14 N_XCSA/LV2_C[4]_XCSA/X_LV2_HA2/M14_d
+ N_XCSA/X_LV2_HA2/N001_XCSA/X_LV2_HA2/M14_g N_GND_XCSA/X_LV2_HA2/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa55/Xao2/M38 N_XADDER/XA55/XAO2/N008_XADDER/Xa55/Xao2/M38_d
+ N_XADDER/GG5_XADDER/Xa55/Xao2/M38_g N_GND_XADDER/Xa55/Xao2/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA0/M18 N_XCSA/X_LV3_FA0/N004_XCSA/X_LV3_FA0/M18_d
+ N_CACC[1]_XCSA/X_LV3_FA0/M18_g N_GND_XCSA/X_LV3_FA0/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA0/M22 N_XCSA/X_LV3_FA0/_SUM_XCSA/X_LV3_FA0/M22_d
+ N_CACC[1]_XCSA/X_LV3_FA0/M22_g N_XCSA/X_LV3_FA0/P005_XCSA/X_LV3_FA0/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV3_FA0/M15 N_XCSA/X_LV3_FA0/_COUT_XCSA/X_LV3_FA0/M15_d
+ N_CACC[1]_XCSA/X_LV3_FA0/M15_g N_XCSA/X_LV3_FA0/N003_XCSA/X_LV3_FA0/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXBOOTH/Xsel21/M3 N_XBOOTH/XSEL21/N002_XBOOTH/Xsel21/M3_d
+ N_XBOOTH/S2_XBOOTH/Xsel21/M3_g N_noxref_2137_XBOOTH/Xsel21/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel11/M3 N_XBOOTH/XSEL11/N002_XBOOTH/Xsel11/M3_d
+ N_XBOOTH/S1_XBOOTH/Xsel11/M3_g N_noxref_2138_XBOOTH/Xsel11/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel01/M3 N_XBOOTH/XSEL01/N002_XBOOTH/Xsel01/M3_d
+ N_XBOOTH/S0_XBOOTH/Xsel01/M3_g N_noxref_2139_XBOOTH/Xsel01/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXADDER/Xa15/Xyb1/Xand1/M16 N_XADDER/PP5_XADDER/Xa15/Xyb1/Xand1/M16_d
+ N_XADDER/XA15/XYB1/N003_XADDER/Xa15/Xyb1/Xand1/M16_g
+ N_GND_XADDER/Xa15/Xyb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd25/M8 N_X02/XD25/N3_X02/xd25/M8_d N_CLK_X02/xd25/M8_g
+ N_X02/XD25/P003_X02/xd25/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa05/Xrb2/M3 N_XADDER/P4_XADDER/Xa05/Xrb2/M3_d
+ N_XADDER/XA05/XRB2/N002_XADDER/Xa05/Xrb2/M3_g N_GND_XADDER/Xa05/Xrb2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xdffb1/M3 N_XBOOTH/XDFFB1/N0_XBOOTH/Xdffb1/M3_d
+ N_B[1]_XBOOTH/Xdffb1/M3_g N_GND_XBOOTH/Xdffb1/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA0/M20 N_XCSA/X_LV3_FA0/N004_XCSA/X_LV3_FA0/M20_d
+ N_PP0[1]_XCSA/X_LV3_FA0/M20_g N_GND_XCSA/X_LV3_FA0/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA0/M23 N_XCSA/X_LV3_FA0/P005_XCSA/X_LV3_FA0/M23_d
+ N_PP0[1]_XCSA/X_LV3_FA0/M23_g N_XCSA/X_LV3_FA0/P006_XCSA/X_LV3_FA0/M23_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA0/M13 N_XCSA/X_LV3_FA0/_COUT_XCSA/X_LV3_FA0/M13_d
+ N_PP0[1]_XCSA/X_LV3_FA0/M13_g N_XCSA/X_LV3_FA0/P004_XCSA/X_LV3_FA0/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA0/M17 N_XCSA/X_LV3_FA0/N003_XCSA/X_LV3_FA0/M17_d
+ N_PP0[1]_XCSA/X_LV3_FA0/M17_g N_GND_XCSA/X_LV3_FA0/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXBOOTH/Xsel21/M4 N_noxref_2137_XBOOTH/Xsel21/M4_d
+ N_XBOOTH/B_D[1]_XBOOTH/Xsel21/M4_g N_GND_XBOOTH/Xsel21/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel11/M4 N_noxref_2138_XBOOTH/Xsel11/M4_d
+ N_XBOOTH/B_D[1]_XBOOTH/Xsel11/M4_g N_GND_XBOOTH/Xsel11/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel01/M4 N_noxref_2139_XBOOTH/Xsel01/M4_d
+ N_XBOOTH/B_D[1]_XBOOTH/Xsel01/M4_g N_GND_XBOOTH/Xsel01/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mX02/xd25/M9 N_X02/XD25/P003_X02/xd25/M9_d N_X02/XD25/N1_X02/xd25/M9_g
+ N_GND_X02/xd25/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.76e-13 PD=2.8e-07 PS=8e-07
mXCSA/Xdffa1/M8 N_XCSA/XDFFA1/N3_XCSA/Xdffa1/M8_d N_CLK_XCSA/Xdffa1/M8_g
+ N_XCSA/XDFFA1/P003_XCSA/Xdffa1/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa14/M8 N_XCSA/XDFFA14/N3_XCSA/Xdffa14/M8_d N_CLK_XCSA/Xdffa14/M8_g
+ N_XCSA/XDFFA14/P003_XCSA/Xdffa14/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xdffb1/M6 N_XBOOTH/XDFFB1/P002_XBOOTH/Xdffb1/M6_d
+ N_CLK_XBOOTH/Xdffb1/M6_g N_GND_XBOOTH/Xdffb1/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXADDER/Xa55/Xao2/Xor1/M16 N_XADDER/GX5[0]_XADDER/Xa55/Xao2/Xor1/M16_d
+ N_XADDER/XA55/XAO2/N008_XADDER/Xa55/Xao2/Xor1/M16_g
+ N_GND_XADDER/Xa55/Xao2/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA0/M19 N_XCSA/X_LV3_FA0/N004_XCSA/X_LV3_FA0/M19_d
+ N_XCSA/LV2_C[1]_XCSA/X_LV3_FA0/M19_g N_GND_XCSA/X_LV3_FA0/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA0/M24 N_XCSA/X_LV3_FA0/P006_XCSA/X_LV3_FA0/M24_d
+ N_XCSA/LV2_C[1]_XCSA/X_LV3_FA0/M24_g N_GND_XCSA/X_LV3_FA0/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA0/M14 N_XCSA/X_LV3_FA0/P004_XCSA/X_LV3_FA0/M14_d
+ N_XCSA/LV2_C[1]_XCSA/X_LV3_FA0/M14_g N_GND_XCSA/X_LV3_FA0/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA0/M16 N_XCSA/X_LV3_FA0/N003_XCSA/X_LV3_FA0/M16_d
+ N_XCSA/LV2_C[1]_XCSA/X_LV3_FA0/M16_g N_GND_XCSA/X_LV3_FA0/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel21/M5 N_XBOOTH/XSEL21/B_XBOOTH/Xsel21/M5_d
+ N_XBOOTH/XSEL21/N002_XBOOTH/Xsel21/M5_g N_GND_XBOOTH/Xsel21/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel11/M5 N_XBOOTH/XSEL11/B_XBOOTH/Xsel11/M5_d
+ N_XBOOTH/XSEL11/N002_XBOOTH/Xsel11/M5_g N_GND_XBOOTH/Xsel11/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel01/M5 N_XBOOTH/XSEL01/B_XBOOTH/Xsel01/M5_d
+ N_XBOOTH/XSEL01/N002_XBOOTH/Xsel01/M5_g N_GND_XBOOTH/Xsel01/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa1/M9 N_XCSA/XDFFA1/P003_XCSA/Xdffa1/M9_d
+ N_XCSA/XDFFA1/N1_XCSA/Xdffa1/M9_g N_GND_XCSA/Xdffa1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/Xdffa14/M9 N_XCSA/XDFFA14/P003_XCSA/Xdffa14/M9_d
+ N_XCSA/XDFFA14/N1_XCSA/Xdffa14/M9_g N_GND_XCSA/Xdffa14/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXADDER/Xa15/Xyb1/M9 N_XADDER/XA15/XYB1/N003_XADDER/Xa15/Xyb1/M9_d
+ N_XADDER/P4_XADDER/Xa15/Xyb1/M9_g
+ N_XADDER/XA15/XYB1/N004_XADDER/Xa15/Xyb1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=9.24e-14 PD=1.44e-06 PS=4.2e-07
mXBOOTH/Xdffb1/M5 N_XBOOTH/XDFFB1/N1_XBOOTH/Xdffb1/M5_d
+ N_XBOOTH/XDFFB1/N0_XBOOTH/Xdffb1/M5_g N_XBOOTH/XDFFB1/P002_XBOOTH/Xdffb1/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV1_FA0/M19 N_XCSA/X_LV1_FA0/N004_XCSA/X_LV1_FA0/M19_d
+ N_PP0[4]_XCSA/X_LV1_FA0/M19_g N_GND_XCSA/X_LV1_FA0/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA0/M24 N_XCSA/X_LV1_FA0/P006_XCSA/X_LV1_FA0/M24_d
+ N_PP0[4]_XCSA/X_LV1_FA0/M24_g N_GND_XCSA/X_LV1_FA0/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA0/M14 N_XCSA/X_LV1_FA0/P004_XCSA/X_LV1_FA0/M14_d
+ N_PP0[4]_XCSA/X_LV1_FA0/M14_g N_GND_XCSA/X_LV1_FA0/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA0/M16 N_XCSA/X_LV1_FA0/N003_XCSA/X_LV1_FA0/M16_d
+ N_PP0[4]_XCSA/X_LV1_FA0/M16_g N_GND_XCSA/X_LV1_FA0/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd25/M11 N_OUT[4]_X02/xd25/M11_d N_X02/XD25/N3_X02/xd25/M11_g
+ N_GND_X02/xd25/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXADDER/Xa05/Xrb2/M1 N_XADDER/XA05/XRB2/N002_XADDER/Xa05/Xrb2/M1_d
+ N_C[4]_XADDER/Xa05/Xrb2/M1_g N_S[4]_XADDER/Xa05/Xrb2/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_FA0/M16 N_XCSA/X_LV2_FA0/N003_XCSA/X_LV2_FA0/M16_d
+ N_XCSA/LV1_C[4]_XCSA/X_LV2_FA0/M16_g N_GND_XCSA/X_LV2_FA0/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV2_FA0/M14 N_XCSA/X_LV2_FA0/P004_XCSA/X_LV2_FA0/M14_d
+ N_XCSA/LV1_C[4]_XCSA/X_LV2_FA0/M14_g N_GND_XCSA/X_LV2_FA0/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_FA0/M24 N_XCSA/X_LV2_FA0/P006_XCSA/X_LV2_FA0/M24_d
+ N_XCSA/LV1_C[4]_XCSA/X_LV2_FA0/M24_g N_GND_XCSA/X_LV2_FA0/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_FA0/M19 N_XCSA/X_LV2_FA0/N004_XCSA/X_LV2_FA0/M19_d
+ N_XCSA/LV1_C[4]_XCSA/X_LV2_FA0/M19_g N_GND_XCSA/X_LV2_FA0/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa15/Xyb1/M10 N_XADDER/XA15/XYB1/N004_XADDER/Xa15/Xyb1/M10_d
+ N_XADDER/P5_XADDER/Xa15/Xyb1/M10_g N_GND_XADDER/Xa15/Xyb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=9.24e-14 AS=2.244e-13
+ PD=4.2e-07 PS=1.46e-06
mXCSA/Xdffa1/M11 N_C[2]_XCSA/Xdffa1/M11_d N_XCSA/XDFFA1/N3_XCSA/Xdffa1/M11_g
+ N_GND_XCSA/Xdffa1/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/Xdffa14/M11 N_S[2]_XCSA/Xdffa14/M11_d N_XCSA/XDFFA14/N3_XCSA/Xdffa14/M11_g
+ N_GND_XCSA/Xdffa14/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/X_LV1_FA0/M20 N_XCSA/X_LV1_FA0/N004_XCSA/X_LV1_FA0/M20_d
+ N_PP1[2]_XCSA/X_LV1_FA0/M20_g N_GND_XCSA/X_LV1_FA0/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV1_FA0/M23 N_XCSA/X_LV1_FA0/P005_XCSA/X_LV1_FA0/M23_d
+ N_PP1[2]_XCSA/X_LV1_FA0/M23_g N_XCSA/X_LV1_FA0/P006_XCSA/X_LV1_FA0/M23_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA0/M13 N_XCSA/X_LV1_FA0/_COUT_XCSA/X_LV1_FA0/M13_d
+ N_PP1[2]_XCSA/X_LV1_FA0/M13_g N_XCSA/X_LV1_FA0/P004_XCSA/X_LV1_FA0/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA0/M17 N_XCSA/X_LV1_FA0/N003_XCSA/X_LV1_FA0/M17_d
+ N_PP1[2]_XCSA/X_LV1_FA0/M17_g N_GND_XCSA/X_LV1_FA0/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXADDER/Xa05/Xrb2/M2 N_XADDER/XA05/XRB2/N002_XADDER/Xa05/Xrb2/M2_d
+ N_S[4]_XADDER/Xa05/Xrb2/M2_g N_C[4]_XADDER/Xa05/Xrb2/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_FA0/M17 N_XCSA/X_LV2_FA0/N003_XCSA/X_LV2_FA0/M17_d
+ N_XCSA/LV1_S[4]_XCSA/X_LV2_FA0/M17_g N_GND_XCSA/X_LV2_FA0/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV2_FA0/M13 N_XCSA/X_LV2_FA0/_COUT_XCSA/X_LV2_FA0/M13_d
+ N_XCSA/LV1_S[4]_XCSA/X_LV2_FA0/M13_g
+ N_XCSA/X_LV2_FA0/P004_XCSA/X_LV2_FA0/M13_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV2_FA0/M23 N_XCSA/X_LV2_FA0/P005_XCSA/X_LV2_FA0/M23_d
+ N_XCSA/LV1_S[4]_XCSA/X_LV2_FA0/M23_g
+ N_XCSA/X_LV2_FA0/P006_XCSA/X_LV2_FA0/M23_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV2_FA0/M20 N_XCSA/X_LV2_FA0/N004_XCSA/X_LV2_FA0/M20_d
+ N_XCSA/LV1_S[4]_XCSA/X_LV2_FA0/M20_g N_GND_XCSA/X_LV2_FA0/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXADDER/Xa64/Xao1/M9 N_XADDER/XA64/XAO1/N003_XADDER/Xa64/Xao1/M9_d
+ N_XADDER/GGG3_XADDER/Xa64/Xao1/M9_g
+ N_XADDER/XA64/XAO1/N004_XADDER/Xa64/Xao1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14 PD=1.44e-06 PS=2.8e-07
mXBOOTH/Xdffb1/M8 N_XBOOTH/XDFFB1/N3_XBOOTH/Xdffb1/M8_d N_CLK_XBOOTH/Xdffb1/M8_g
+ N_XBOOTH/XDFFB1/P003_XBOOTH/Xdffb1/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mX02/xd26/M3 N_X02/XD26/N0_X02/xd26/M3_d N_OUT1[5]_X02/xd26/M3_g
+ N_GND_X02/xd26/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA0/M18 N_XCSA/X_LV1_FA0/N004_XCSA/X_LV1_FA0/M18_d
+ N_PP2[0]_XCSA/X_LV1_FA0/M18_g N_GND_XCSA/X_LV1_FA0/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV1_FA0/M22 N_XCSA/X_LV1_FA0/_SUM_XCSA/X_LV1_FA0/M22_d
+ N_PP2[0]_XCSA/X_LV1_FA0/M22_g N_XCSA/X_LV1_FA0/P005_XCSA/X_LV1_FA0/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV1_FA0/M15 N_XCSA/X_LV1_FA0/_COUT_XCSA/X_LV1_FA0/M15_d
+ N_PP2[0]_XCSA/X_LV1_FA0/M15_g N_XCSA/X_LV1_FA0/N003_XCSA/X_LV1_FA0/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXADDER/Xa64/Xao1/M10 N_XADDER/XA64/XAO1/N004_XADDER/Xa64/Xao1/M10_d
+ N_XADDER/P4_XADDER/Xa64/Xao1/M10_g N_GND_XADDER/Xa64/Xao1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.86e-13
+ PD=2.8e-07 PS=1.74e-06
mXCSA/X_LV2_FA0/M15 N_XCSA/X_LV2_FA0/_COUT_XCSA/X_LV2_FA0/M15_d
+ N_A_D[5]_XCSA/X_LV2_FA0/M15_g N_XCSA/X_LV2_FA0/N003_XCSA/X_LV2_FA0/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV2_FA0/M22 N_XCSA/X_LV2_FA0/_SUM_XCSA/X_LV2_FA0/M22_d
+ N_A_D[5]_XCSA/X_LV2_FA0/M22_g N_XCSA/X_LV2_FA0/P005_XCSA/X_LV2_FA0/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV2_FA0/M18 N_XCSA/X_LV2_FA0/N004_XCSA/X_LV2_FA0/M18_d
+ N_A_D[5]_XCSA/X_LV2_FA0/M18_g N_GND_XCSA/X_LV2_FA0/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXBOOTH/Xsel21/M12 N_XBOOTH/XSEL21/N004_XBOOTH/Xsel21/M12_d
+ N_A_D[5]_XBOOTH/Xsel21/M12_g N_XBOOTH/XSEL21/B_XBOOTH/Xsel21/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel11/M12 N_XBOOTH/XSEL11/N004_XBOOTH/Xsel11/M12_d
+ N_A_D[3]_XBOOTH/Xsel11/M12_g N_XBOOTH/XSEL11/B_XBOOTH/Xsel11/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel01/M12 N_XBOOTH/XSEL01/N004_XBOOTH/Xsel01/M12_d
+ N_A_D[1]_XBOOTH/Xsel01/M12_g N_XBOOTH/XSEL01/B_XBOOTH/Xsel01/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_HA1/M11 N_XCSA/X_LV3_HA1/P001_XCSA/X_LV3_HA1/M11_d
+ N_XCSA/LV2_S[2]_XCSA/X_LV3_HA1/M11_g N_GND_XCSA/X_LV3_HA1/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV3_HA1/X_xor/M2 N_XCSA/X_LV3_HA1/X_XOR/N002_XCSA/X_LV3_HA1/X_xor/M2_d
+ N_XCSA/LV2_S[2]_XCSA/X_LV3_HA1/X_xor/M2_g N_CACC[2]_XCSA/X_LV3_HA1/X_xor/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXBOOTH/Xdffb1/M9 N_XBOOTH/XDFFB1/P003_XBOOTH/Xdffb1/M9_d
+ N_XBOOTH/XDFFB1/N1_XBOOTH/Xdffb1/M9_g N_GND_XBOOTH/Xdffb1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXADDER/Xa15/Xyb2/M10 N_XADDER/XA15/XYB2/N004_XADDER/Xa15/Xyb2/M10_d
+ N_XADDER/P5_XADDER/Xa15/Xyb2/M10_g N_GND_XADDER/Xa15/Xyb2/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXCSA/Xdffa2/M3 N_XCSA/XDFFA2/N0_XCSA/Xdffa2/M3_d
+ N_XCSA/LV3_C[3]_XCSA/Xdffa2/M3_g N_GND_XCSA/Xdffa2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa15/M3 N_XCSA/XDFFA15/N0_XCSA/Xdffa15/M3_d
+ N_XCSA/LV3_S[3]_XCSA/Xdffa15/M3_g N_GND_XCSA/Xdffa15/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd26/M6 N_X02/XD26/P002_X02/xd26/M6_d N_CLK_X02/xd26/M6_g
+ N_GND_X02/xd26/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/X_LV1_FA0/M21 N_XCSA/X_LV1_FA0/_SUM_XCSA/X_LV1_FA0/M21_d
+ N_XCSA/X_LV1_FA0/_COUT_XCSA/X_LV1_FA0/M21_g
+ N_XCSA/X_LV1_FA0/N004_XCSA/X_LV1_FA0/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXADDER/Xa15/Xyb2/M9 N_XADDER/XA15/XYB2/N003_XADDER/Xa15/Xyb2/M9_d
+ N_XADDER/G4_XADDER/Xa15/Xyb2/M9_g
+ N_XADDER/XA15/XYB2/N004_XADDER/Xa15/Xyb2/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=6.16e-14 PD=1.74e-06 PS=2.8e-07
mXBOOTH/Xsel21/M11 N_XBOOTH/XSEL21/N004_XBOOTH/Xsel21/M11_d
+ N_XBOOTH/XSEL21/B_XBOOTH/Xsel21/M11_g N_A_D[5]_XBOOTH/Xsel21/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel11/M11 N_XBOOTH/XSEL11/N004_XBOOTH/Xsel11/M11_d
+ N_XBOOTH/XSEL11/B_XBOOTH/Xsel11/M11_g N_A_D[3]_XBOOTH/Xsel11/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel01/M11 N_XBOOTH/XSEL01/N004_XBOOTH/Xsel01/M11_d
+ N_XBOOTH/XSEL01/B_XBOOTH/Xsel01/M11_g N_A_D[1]_XBOOTH/Xsel01/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_HA1/M12 N_XCSA/X_LV3_HA1/N001_XCSA/X_LV3_HA1/M12_d
+ N_CACC[2]_XCSA/X_LV3_HA1/M12_g N_XCSA/X_LV3_HA1/P001_XCSA/X_LV3_HA1/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_HA1/X_xor/M1 N_XCSA/X_LV3_HA1/X_XOR/N002_XCSA/X_LV3_HA1/X_xor/M1_d
+ N_CACC[2]_XCSA/X_LV3_HA1/X_xor/M1_g N_XCSA/LV2_S[2]_XCSA/X_LV3_HA1/X_xor/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa05/Xrb1/M10 N_XADDER/XA05/XRB1/N004_XADDER/Xa05/Xrb1/M10_d
+ N_S[4]_XADDER/Xa05/Xrb1/M10_g N_GND_XADDER/Xa05/Xrb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXCSA/X_LV2_FA0/M21 N_XCSA/X_LV2_FA0/_SUM_XCSA/X_LV2_FA0/M21_d
+ N_XCSA/X_LV2_FA0/_COUT_XCSA/X_LV2_FA0/M21_g
+ N_XCSA/X_LV2_FA0/N004_XCSA/X_LV2_FA0/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mX02/xd26/M5 N_X02/XD26/N1_X02/xd26/M5_d N_X02/XD26/N0_X02/xd26/M5_g
+ N_X02/XD26/P002_X02/xd26/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xdffb1/M11 N_XBOOTH/B_D[1]_XBOOTH/Xdffb1/M11_d
+ N_XBOOTH/XDFFB1/N3_XBOOTH/Xdffb1/M11_g N_GND_XBOOTH/Xdffb1/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXADDER/Xa75/M3 N_OUT1[5]_XADDER/Xa75/M3_d N_XADDER/XA75/N002_XADDER/Xa75/M3_g
+ N_GND_XADDER/Xa75/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa2/M6 N_XCSA/XDFFA2/P002_XCSA/Xdffa2/M6_d N_CLK_XCSA/Xdffa2/M6_g
+ N_GND_XCSA/Xdffa2/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/Xdffa15/M6 N_XCSA/XDFFA15/P002_XCSA/Xdffa15/M6_d N_CLK_XCSA/Xdffa15/M6_g
+ N_GND_XCSA/Xdffa15/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXADDER/Xa05/Xrb1/M9 N_XADDER/XA05/XRB1/N003_XADDER/Xa05/Xrb1/M9_d
+ N_C[4]_XADDER/Xa05/Xrb1/M9_g N_XADDER/XA05/XRB1/N004_XADDER/Xa05/Xrb1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14
+ PD=1.44e-06 PS=2.8e-07
mXCSA/X_LV1_FA0/M26 N_XCSA/LV1_C[5]_XCSA/X_LV1_FA0/M26_d
+ N_XCSA/X_LV1_FA0/_COUT_XCSA/X_LV1_FA0/M26_g N_GND_XCSA/X_LV1_FA0/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_FA0/M26 N_XCSA/LV2_C[5]_XCSA/X_LV2_FA0/M26_d
+ N_XCSA/X_LV2_FA0/_COUT_XCSA/X_LV2_FA0/M26_g N_GND_XCSA/X_LV2_FA0/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa64/Xao1/Xand1/M16 N_XADDER/XA64/OUT1_XADDER/Xa64/Xao1/Xand1/M16_d
+ N_XADDER/XA64/XAO1/N003_XADDER/Xa64/Xao1/Xand1/M16_g
+ N_GND_XADDER/Xa64/Xao1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa2/M5 N_XCSA/XDFFA2/N1_XCSA/Xdffa2/M5_d
+ N_XCSA/XDFFA2/N0_XCSA/Xdffa2/M5_g N_XCSA/XDFFA2/P002_XCSA/Xdffa2/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa15/M5 N_XCSA/XDFFA15/N1_XCSA/Xdffa15/M5_d
+ N_XCSA/XDFFA15/N0_XCSA/Xdffa15/M5_g N_XCSA/XDFFA15/P002_XCSA/Xdffa15/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel21/M13 N_PP2[1]_XBOOTH/Xsel21/M13_d
+ N_XBOOTH/XSEL21/N004_XBOOTH/Xsel21/M13_g N_GND_XBOOTH/Xsel21/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel11/M13 N_PP1[1]_XBOOTH/Xsel11/M13_d
+ N_XBOOTH/XSEL11/N004_XBOOTH/Xsel11/M13_g N_GND_XBOOTH/Xsel11/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel01/M13 N_PP0[1]_XBOOTH/Xsel01/M13_d
+ N_XBOOTH/XSEL01/N004_XBOOTH/Xsel01/M13_g N_GND_XBOOTH/Xsel01/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA0/M25 N_XCSA/LV1_S[4]_XCSA/X_LV1_FA0/M25_d
+ N_XCSA/X_LV1_FA0/_SUM_XCSA/X_LV1_FA0/M25_g N_GND_XCSA/X_LV1_FA0/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_HA1/M14 N_XCSA/LV3_C[3]_XCSA/X_LV3_HA1/M14_d
+ N_XCSA/X_LV3_HA1/N001_XCSA/X_LV3_HA1/M14_g N_GND_XCSA/X_LV3_HA1/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_HA1/X_xor/M3 N_XCSA/LV3_S[2]_XCSA/X_LV3_HA1/X_xor/M3_d
+ N_XCSA/X_LV3_HA1/X_XOR/N002_XCSA/X_LV3_HA1/X_xor/M3_g
+ N_GND_XCSA/X_LV3_HA1/X_xor/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_FA0/M25 N_XCSA/LV2_S[4]_XCSA/X_LV2_FA0/M25_d
+ N_XCSA/X_LV2_FA0/_SUM_XCSA/X_LV2_FA0/M25_g N_GND_XCSA/X_LV2_FA0/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa15/Xyb2/Xand1/M16 N_XADDER/XA15/T1_XADDER/Xa15/Xyb2/Xand1/M16_d
+ N_XADDER/XA15/XYB2/N003_XADDER/Xa15/Xyb2/Xand1/M16_g
+ N_GND_XADDER/Xa15/Xyb2/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd26/M8 N_X02/XD26/N3_X02/xd26/M8_d N_CLK_X02/xd26/M8_g
+ N_X02/XD26/P003_X02/xd26/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa05/Xrb1/Xand1/M16 N_XADDER/G4_XADDER/Xa05/Xrb1/Xand1/M16_d
+ N_XADDER/XA05/XRB1/N003_XADDER/Xa05/Xrb1/Xand1/M16_g
+ N_GND_XADDER/Xa05/Xrb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd26/M9 N_X02/XD26/P003_X02/xd26/M9_d N_X02/XD26/N1_X02/xd26/M9_g
+ N_GND_X02/xd26/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.76e-13 PD=2.8e-07 PS=8e-07
mXADDER/Xa64/Xao2/M37 N_XADDER/XA64/XAO2/N008_XADDER/Xa64/Xao2/M37_d
+ N_XADDER/XA64/OUT1_XADDER/Xa64/Xao2/M37_g N_GND_XADDER/Xa64/Xao2/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa2/M8 N_XCSA/XDFFA2/N3_XCSA/Xdffa2/M8_d N_CLK_XCSA/Xdffa2/M8_g
+ N_XCSA/XDFFA2/P003_XCSA/Xdffa2/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa15/M8 N_XCSA/XDFFA15/N3_XCSA/Xdffa15/M8_d N_CLK_XCSA/Xdffa15/M8_g
+ N_XCSA/XDFFA15/P003_XCSA/Xdffa15/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa75/M1 N_XADDER/XA75/N002_XADDER/Xa75/M1_d N_XADDER/P5_XADDER/Xa75/M1_g
+ N_XADDER/GX6[1]_XADDER/Xa75/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=2.332e-13 PD=5.4e-07 PS=1.5e-06
mXCSA/Xdffa2/M9 N_XCSA/XDFFA2/P003_XCSA/Xdffa2/M9_d
+ N_XCSA/XDFFA2/N1_XCSA/Xdffa2/M9_g N_GND_XCSA/Xdffa2/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/Xdffa15/M9 N_XCSA/XDFFA15/P003_XCSA/Xdffa15/M9_d
+ N_XCSA/XDFFA15/N1_XCSA/Xdffa15/M9_g N_GND_XCSA/Xdffa15/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXADDER/Xa64/Xao2/M38 N_XADDER/XA64/XAO2/N008_XADDER/Xa64/Xao2/M38_d
+ N_XADDER/G4_XADDER/Xa64/Xao2/M38_g N_GND_XADDER/Xa64/Xao2/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa15/Xyb3/M37 N_XADDER/XA15/XYB3/N008_XADDER/Xa15/Xyb3/M37_d
+ N_XADDER/XA15/T1_XADDER/Xa15/Xyb3/M37_g N_GND_XADDER/Xa15/Xyb3/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa75/M2 N_XADDER/XA75/N002_XADDER/Xa75/M2_d
+ N_XADDER/GX6[1]_XADDER/Xa75/M2_g N_XADDER/P5_XADDER/Xa75/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mX02/xd26/M11 N_OUT[5]_X02/xd26/M11_d N_X02/XD26/N3_X02/xd26/M11_g
+ N_GND_X02/xd26/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXBOOTH/Xsel22/M2 N_noxref_2164_XBOOTH/Xsel22/M2_d
+ N_XBOOTH/B_D[1]_XBOOTH/Xsel22/M2_g N_GND_XBOOTH/Xsel22/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel12/M2 N_noxref_2165_XBOOTH/Xsel12/M2_d
+ N_XBOOTH/B_D[1]_XBOOTH/Xsel12/M2_g N_GND_XBOOTH/Xsel12/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel02/M2 N_noxref_2166_XBOOTH/Xsel02/M2_d
+ N_XBOOTH/B_D[1]_XBOOTH/Xsel02/M2_g N_GND_XBOOTH/Xsel02/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_HA3/X_xor/M2 N_XCSA/X_LV2_HA3/X_XOR/N002_XCSA/X_LV2_HA3/X_xor/M2_d
+ N_XCSA/LV1_C[5]_XCSA/X_LV2_HA3/X_xor/M2_g
+ N_XCSA/LV1_S[5]_XCSA/X_LV2_HA3/X_xor/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13 PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA3/M11 N_XCSA/X_LV2_HA3/P001_XCSA/X_LV2_HA3/M11_d
+ N_XCSA/LV1_C[5]_XCSA/X_LV2_HA3/M11_g N_GND_XCSA/X_LV2_HA3/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV3_FA1/M25 N_XCSA/LV3_S[3]_XCSA/X_LV3_FA1/M25_d
+ N_XCSA/X_LV3_FA1/_SUM_XCSA/X_LV3_FA1/M25_g N_GND_XCSA/X_LV3_FA1/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA1/M19 N_XCSA/X_LV1_FA1/N004_XCSA/X_LV1_FA1/M19_d
+ N_PP0[5]_XCSA/X_LV1_FA1/M19_g N_GND_XCSA/X_LV1_FA1/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA1/M24 N_XCSA/X_LV1_FA1/P006_XCSA/X_LV1_FA1/M24_d
+ N_PP0[5]_XCSA/X_LV1_FA1/M24_g N_GND_XCSA/X_LV1_FA1/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA1/M14 N_XCSA/X_LV1_FA1/P004_XCSA/X_LV1_FA1/M14_d
+ N_PP0[5]_XCSA/X_LV1_FA1/M14_g N_GND_XCSA/X_LV1_FA1/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA1/M16 N_XCSA/X_LV1_FA1/N003_XCSA/X_LV1_FA1/M16_d
+ N_PP0[5]_XCSA/X_LV1_FA1/M16_g N_GND_XCSA/X_LV1_FA1/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa06/Xrb2/M3 N_XADDER/P5_XADDER/Xa06/Xrb2/M3_d
+ N_XADDER/XA06/XRB2/N002_XADDER/Xa06/Xrb2/M3_g N_GND_XADDER/Xa06/Xrb2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa15/Xyb3/M38 N_XADDER/XA15/XYB3/N008_XADDER/Xa15/Xyb3/M38_d
+ N_XADDER/G5_XADDER/Xa15/Xyb3/M38_g N_GND_XADDER/Xa15/Xyb3/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa2/M11 N_C[3]_XCSA/Xdffa2/M11_d N_XCSA/XDFFA2/N3_XCSA/Xdffa2/M11_g
+ N_GND_XCSA/Xdffa2/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/Xdffa15/M11 N_S[3]_XCSA/Xdffa15/M11_d N_XCSA/XDFFA15/N3_XCSA/Xdffa15/M11_g
+ N_GND_XCSA/Xdffa15/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXBOOTH/Xsel22/M1 N_XBOOTH/XSEL22/N002_XBOOTH/Xsel22/M1_d
+ N_XBOOTH/D2_XBOOTH/Xsel22/M1_g N_noxref_2164_XBOOTH/Xsel22/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel12/M1 N_XBOOTH/XSEL12/N002_XBOOTH/Xsel12/M1_d
+ N_XBOOTH/D1_XBOOTH/Xsel12/M1_g N_noxref_2165_XBOOTH/Xsel12/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel02/M1 N_XBOOTH/XSEL02/N002_XBOOTH/Xsel02/M1_d
+ N_XBOOTH/D0_XBOOTH/Xsel02/M1_g N_noxref_2166_XBOOTH/Xsel02/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXCSA/X_LV2_HA3/X_xor/M1 N_XCSA/X_LV2_HA3/X_XOR/N002_XCSA/X_LV2_HA3/X_xor/M1_d
+ N_XCSA/LV1_S[5]_XCSA/X_LV2_HA3/X_xor/M1_g
+ N_XCSA/LV1_C[5]_XCSA/X_LV2_HA3/X_xor/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_HA3/M12 N_XCSA/X_LV2_HA3/N001_XCSA/X_LV2_HA3/M12_d
+ N_XCSA/LV1_S[5]_XCSA/X_LV2_HA3/M12_g
+ N_XCSA/X_LV2_HA3/P001_XCSA/X_LV2_HA3/M12_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA1/M26 N_XCSA/LV3_C[4]_XCSA/X_LV3_FA1/M26_d
+ N_XCSA/X_LV3_FA1/_COUT_XCSA/X_LV3_FA1/M26_g N_GND_XCSA/X_LV3_FA1/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA1/M20 N_XCSA/X_LV1_FA1/N004_XCSA/X_LV1_FA1/M20_d
+ N_PP1[3]_XCSA/X_LV1_FA1/M20_g N_GND_XCSA/X_LV1_FA1/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV1_FA1/M23 N_XCSA/X_LV1_FA1/P005_XCSA/X_LV1_FA1/M23_d
+ N_PP1[3]_XCSA/X_LV1_FA1/M23_g N_XCSA/X_LV1_FA1/P006_XCSA/X_LV1_FA1/M23_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA1/M13 N_XCSA/X_LV1_FA1/_COUT_XCSA/X_LV1_FA1/M13_d
+ N_PP1[3]_XCSA/X_LV1_FA1/M13_g N_XCSA/X_LV1_FA1/P004_XCSA/X_LV1_FA1/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA1/M17 N_XCSA/X_LV1_FA1/N003_XCSA/X_LV1_FA1/M17_d
+ N_PP1[3]_XCSA/X_LV1_FA1/M17_g N_GND_XCSA/X_LV1_FA1/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXADDER/Xa64/Xao2/Xor1/M16 N_XADDER/GX6[1]_XADDER/Xa64/Xao2/Xor1/M16_d
+ N_XADDER/XA64/XAO2/N008_XADDER/Xa64/Xao2/Xor1/M16_g
+ N_GND_XADDER/Xa64/Xao2/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd27/M3 N_X02/XD27/N0_X02/xd27/M3_d N_OUT1[6]_X02/xd27/M3_g
+ N_GND_X02/xd27/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel22/M3 N_XBOOTH/XSEL22/N002_XBOOTH/Xsel22/M3_d
+ N_XBOOTH/S2_XBOOTH/Xsel22/M3_g N_noxref_2171_XBOOTH/Xsel22/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel12/M3 N_XBOOTH/XSEL12/N002_XBOOTH/Xsel12/M3_d
+ N_XBOOTH/S1_XBOOTH/Xsel12/M3_g N_noxref_2172_XBOOTH/Xsel12/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel02/M3 N_XBOOTH/XSEL02/N002_XBOOTH/Xsel02/M3_d
+ N_XBOOTH/S0_XBOOTH/Xsel02/M3_g N_noxref_2173_XBOOTH/Xsel02/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xdffb2/M3 N_XBOOTH/XDFFB2/N0_XBOOTH/Xdffb2/M3_d
+ N_B[2]_XBOOTH/Xdffb2/M3_g N_GND_XBOOTH/Xdffb2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA1/M21 N_XCSA/X_LV3_FA1/_SUM_XCSA/X_LV3_FA1/M21_d
+ N_XCSA/X_LV3_FA1/_COUT_XCSA/X_LV3_FA1/M21_g
+ N_XCSA/X_LV3_FA1/N004_XCSA/X_LV3_FA1/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXCSA/X_LV1_FA1/M18 N_XCSA/X_LV1_FA1/N004_XCSA/X_LV1_FA1/M18_d
+ N_PP2[1]_XCSA/X_LV1_FA1/M18_g N_GND_XCSA/X_LV1_FA1/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV1_FA1/M22 N_XCSA/X_LV1_FA1/_SUM_XCSA/X_LV1_FA1/M22_d
+ N_PP2[1]_XCSA/X_LV1_FA1/M22_g N_XCSA/X_LV1_FA1/P005_XCSA/X_LV1_FA1/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV1_FA1/M15 N_XCSA/X_LV1_FA1/_COUT_XCSA/X_LV1_FA1/M15_d
+ N_PP2[1]_XCSA/X_LV1_FA1/M15_g N_XCSA/X_LV1_FA1/N003_XCSA/X_LV1_FA1/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXADDER/Xa06/Xrb2/M1 N_XADDER/XA06/XRB2/N002_XADDER/Xa06/Xrb2/M1_d
+ N_C[5]_XADDER/Xa06/Xrb2/M1_g N_S[5]_XADDER/Xa06/Xrb2/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa15/Xyb3/Xor1/M16 N_XADDER/GG5_XADDER/Xa15/Xyb3/Xor1/M16_d
+ N_XADDER/XA15/XYB3/N008_XADDER/Xa15/Xyb3/Xor1/M16_g
+ N_GND_XADDER/Xa15/Xyb3/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa3/M3 N_XCSA/XDFFA3/N0_XCSA/Xdffa3/M3_d
+ N_XCSA/LV3_C[4]_XCSA/Xdffa3/M3_g N_GND_XCSA/Xdffa3/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa16/M3 N_XCSA/XDFFA16/N0_XCSA/Xdffa16/M3_d
+ N_XCSA/LV3_S[4]_XCSA/Xdffa16/M3_g N_GND_XCSA/Xdffa16/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa37/Xao1/M9 N_XADDER/XA37/XAO1/N003_XADDER/Xa37/Xao1/M9_d
+ N_XADDER/GGG3_XADDER/Xa37/Xao1/M9_g
+ N_XADDER/XA37/XAO1/N004_XADDER/Xa37/Xao1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14 PD=1.44e-06 PS=2.8e-07
mX02/xd27/M6 N_X02/XD27/P002_X02/xd27/M6_d N_CLK_X02/xd27/M6_g
+ N_GND_X02/xd27/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXBOOTH/Xsel22/M4 N_noxref_2171_XBOOTH/Xsel22/M4_d
+ N_XBOOTH/B_D[2]_XBOOTH/Xsel22/M4_g N_GND_XBOOTH/Xsel22/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel12/M4 N_noxref_2172_XBOOTH/Xsel12/M4_d
+ N_XBOOTH/B_D[2]_XBOOTH/Xsel12/M4_g N_GND_XBOOTH/Xsel12/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel02/M4 N_noxref_2173_XBOOTH/Xsel02/M4_d
+ N_XBOOTH/B_D[2]_XBOOTH/Xsel02/M4_g N_GND_XBOOTH/Xsel02/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xdffb2/M6 N_XBOOTH/XDFFB2/P002_XBOOTH/Xdffb2/M6_d
+ N_CLK_XBOOTH/Xdffb2/M6_g N_GND_XBOOTH/Xdffb2/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXCSA/X_LV2_HA3/X_xor/M3 N_XCSA/LV2_S[5]_XCSA/X_LV2_HA3/X_xor/M3_d
+ N_XCSA/X_LV2_HA3/X_XOR/N002_XCSA/X_LV2_HA3/X_xor/M3_g
+ N_GND_XCSA/X_LV2_HA3/X_xor/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA3/M14 N_XCSA/LV2_C[6]_XCSA/X_LV2_HA3/M14_d
+ N_XCSA/X_LV2_HA3/N001_XCSA/X_LV2_HA3/M14_g N_GND_XCSA/X_LV2_HA3/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA1/M18 N_XCSA/X_LV3_FA1/N004_XCSA/X_LV3_FA1/M18_d
+ N_CACC[3]_XCSA/X_LV3_FA1/M18_g N_GND_XCSA/X_LV3_FA1/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA1/M22 N_XCSA/X_LV3_FA1/_SUM_XCSA/X_LV3_FA1/M22_d
+ N_CACC[3]_XCSA/X_LV3_FA1/M22_g N_XCSA/X_LV3_FA1/P005_XCSA/X_LV3_FA1/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV3_FA1/M15 N_XCSA/X_LV3_FA1/_COUT_XCSA/X_LV3_FA1/M15_d
+ N_CACC[3]_XCSA/X_LV3_FA1/M15_g N_XCSA/X_LV3_FA1/N003_XCSA/X_LV3_FA1/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXADDER/Xa37/Xao1/M10 N_XADDER/XA37/XAO1/N004_XADDER/Xa37/Xao1/M10_d
+ N_XADDER/PPP7_XADDER/Xa37/Xao1/M10_g N_GND_XADDER/Xa37/Xao1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.86e-13
+ PD=2.8e-07 PS=1.74e-06
mX02/xd27/M5 N_X02/XD27/N1_X02/xd27/M5_d N_X02/XD27/N0_X02/xd27/M5_g
+ N_X02/XD27/P002_X02/xd27/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa06/Xrb2/M2 N_XADDER/XA06/XRB2/N002_XADDER/Xa06/Xrb2/M2_d
+ N_S[5]_XADDER/Xa06/Xrb2/M2_g N_C[5]_XADDER/Xa06/Xrb2/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV1_FA1/M21 N_XCSA/X_LV1_FA1/_SUM_XCSA/X_LV1_FA1/M21_d
+ N_XCSA/X_LV1_FA1/_COUT_XCSA/X_LV1_FA1/M21_g
+ N_XCSA/X_LV1_FA1/N004_XCSA/X_LV1_FA1/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXBOOTH/Xdffb2/M5 N_XBOOTH/XDFFB2/N1_XBOOTH/Xdffb2/M5_d
+ N_XBOOTH/XDFFB2/N0_XBOOTH/Xdffb2/M5_g N_XBOOTH/XDFFB2/P002_XBOOTH/Xdffb2/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa3/M6 N_XCSA/XDFFA3/P002_XCSA/Xdffa3/M6_d N_CLK_XCSA/Xdffa3/M6_g
+ N_GND_XCSA/Xdffa3/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/Xdffa16/M6 N_XCSA/XDFFA16/P002_XCSA/Xdffa16/M6_d N_CLK_XCSA/Xdffa16/M6_g
+ N_GND_XCSA/Xdffa16/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXBOOTH/Xsel22/M5 N_XBOOTH/XSEL22/B_XBOOTH/Xsel22/M5_d
+ N_XBOOTH/XSEL22/N002_XBOOTH/Xsel22/M5_g N_GND_XBOOTH/Xsel22/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel12/M5 N_XBOOTH/XSEL12/B_XBOOTH/Xsel12/M5_d
+ N_XBOOTH/XSEL12/N002_XBOOTH/Xsel12/M5_g N_GND_XBOOTH/Xsel12/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel02/M5 N_XBOOTH/XSEL02/B_XBOOTH/Xsel02/M5_d
+ N_XBOOTH/XSEL02/N002_XBOOTH/Xsel02/M5_g N_GND_XBOOTH/Xsel02/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa27/Xyb1/Xand1/M16 N_XADDER/PPP7_XADDER/Xa27/Xyb1/Xand1/M16_d
+ N_XADDER/XA27/XYB1/N003_XADDER/Xa27/Xyb1/Xand1/M16_g
+ N_GND_XADDER/Xa27/Xyb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa3/M5 N_XCSA/XDFFA3/N1_XCSA/Xdffa3/M5_d
+ N_XCSA/XDFFA3/N0_XCSA/Xdffa3/M5_g N_XCSA/XDFFA3/P002_XCSA/Xdffa3/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa16/M5 N_XCSA/XDFFA16/N1_XCSA/Xdffa16/M5_d
+ N_XCSA/XDFFA16/N0_XCSA/Xdffa16/M5_g N_XCSA/XDFFA16/P002_XCSA/Xdffa16/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV3_FA1/M20 N_XCSA/X_LV3_FA1/N004_XCSA/X_LV3_FA1/M20_d
+ N_XCSA/LV2_S[3]_XCSA/X_LV3_FA1/M20_g N_GND_XCSA/X_LV3_FA1/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA1/M23 N_XCSA/X_LV3_FA1/P005_XCSA/X_LV3_FA1/M23_d
+ N_XCSA/LV2_S[3]_XCSA/X_LV3_FA1/M23_g
+ N_XCSA/X_LV3_FA1/P006_XCSA/X_LV3_FA1/M23_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA1/M13 N_XCSA/X_LV3_FA1/_COUT_XCSA/X_LV3_FA1/M13_d
+ N_XCSA/LV2_S[3]_XCSA/X_LV3_FA1/M13_g
+ N_XCSA/X_LV3_FA1/P004_XCSA/X_LV3_FA1/M13_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA1/M17 N_XCSA/X_LV3_FA1/N003_XCSA/X_LV3_FA1/M17_d
+ N_XCSA/LV2_S[3]_XCSA/X_LV3_FA1/M17_g N_GND_XCSA/X_LV3_FA1/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA1/M26 N_XCSA/LV1_C[6]_XCSA/X_LV1_FA1/M26_d
+ N_XCSA/X_LV1_FA1/_COUT_XCSA/X_LV1_FA1/M26_g N_GND_XCSA/X_LV1_FA1/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA1/M19 N_XCSA/X_LV3_FA1/N004_XCSA/X_LV3_FA1/M19_d
+ N_XCSA/LV2_C[3]_XCSA/X_LV3_FA1/M19_g N_GND_XCSA/X_LV3_FA1/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA1/M24 N_XCSA/X_LV3_FA1/P006_XCSA/X_LV3_FA1/M24_d
+ N_XCSA/LV2_C[3]_XCSA/X_LV3_FA1/M24_g N_GND_XCSA/X_LV3_FA1/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA1/M14 N_XCSA/X_LV3_FA1/P004_XCSA/X_LV3_FA1/M14_d
+ N_XCSA/LV2_C[3]_XCSA/X_LV3_FA1/M14_g N_GND_XCSA/X_LV3_FA1/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA1/M16 N_XCSA/X_LV3_FA1/N003_XCSA/X_LV3_FA1/M16_d
+ N_XCSA/LV2_C[3]_XCSA/X_LV3_FA1/M16_g N_GND_XCSA/X_LV3_FA1/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd27/M8 N_X02/XD27/N3_X02/xd27/M8_d N_CLK_X02/xd27/M8_g
+ N_X02/XD27/P003_X02/xd27/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV1_FA1/M25 N_XCSA/LV1_S[5]_XCSA/X_LV1_FA1/M25_d
+ N_XCSA/X_LV1_FA1/_SUM_XCSA/X_LV1_FA1/M25_g N_GND_XCSA/X_LV1_FA1/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xdffb2/M8 N_XBOOTH/XDFFB2/N3_XBOOTH/Xdffb2/M8_d N_CLK_XBOOTH/Xdffb2/M8_g
+ N_XBOOTH/XDFFB2/P003_XBOOTH/Xdffb2/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa37/Xao1/Xand1/M16 N_XADDER/XA37/OUT1_XADDER/Xa37/Xao1/Xand1/M16_d
+ N_XADDER/XA37/XAO1/N003_XADDER/Xa37/Xao1/Xand1/M16_g
+ N_GND_XADDER/Xa37/Xao1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa06/Xrb1/M10 N_XADDER/XA06/XRB1/N004_XADDER/Xa06/Xrb1/M10_d
+ N_S[5]_XADDER/Xa06/Xrb1/M10_g N_GND_XADDER/Xa06/Xrb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXADDER/Xa27/Xyb1/M9 N_XADDER/XA27/XYB1/N003_XADDER/Xa27/Xyb1/M9_d
+ N_XADDER/PP5_XADDER/Xa27/Xyb1/M9_g
+ N_XADDER/XA27/XYB1/N004_XADDER/Xa27/Xyb1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=9.24e-14 PD=1.44e-06 PS=4.2e-07
mX02/xd27/M9 N_X02/XD27/P003_X02/xd27/M9_d N_X02/XD27/N1_X02/xd27/M9_g
+ N_GND_X02/xd27/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.76e-13 PD=2.8e-07 PS=8e-07
mXBOOTH/Xdffb2/M9 N_XBOOTH/XDFFB2/P003_XBOOTH/Xdffb2/M9_d
+ N_XBOOTH/XDFFB2/N1_XBOOTH/Xdffb2/M9_g N_GND_XBOOTH/Xdffb2/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/Xdffa3/M8 N_XCSA/XDFFA3/N3_XCSA/Xdffa3/M8_d N_CLK_XCSA/Xdffa3/M8_g
+ N_XCSA/XDFFA3/P003_XCSA/Xdffa3/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa06/Xrb1/M9 N_XADDER/XA06/XRB1/N003_XADDER/Xa06/Xrb1/M9_d
+ N_C[5]_XADDER/Xa06/Xrb1/M9_g N_XADDER/XA06/XRB1/N004_XADDER/Xa06/Xrb1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14
+ PD=1.44e-06 PS=2.8e-07
mXCSA/Xdffa16/M8 N_XCSA/XDFFA16/N3_XCSA/Xdffa16/M8_d N_CLK_XCSA/Xdffa16/M8_g
+ N_XCSA/XDFFA16/P003_XCSA/Xdffa16/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel22/M12 N_XBOOTH/XSEL22/N004_XBOOTH/Xsel22/M12_d
+ N_A_D[5]_XBOOTH/Xsel22/M12_g N_XBOOTH/XSEL22/B_XBOOTH/Xsel22/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel12/M12 N_XBOOTH/XSEL12/N004_XBOOTH/Xsel12/M12_d
+ N_A_D[3]_XBOOTH/Xsel12/M12_g N_XBOOTH/XSEL12/B_XBOOTH/Xsel12/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel02/M12 N_XBOOTH/XSEL02/N004_XBOOTH/Xsel02/M12_d
+ N_A_D[1]_XBOOTH/Xsel02/M12_g N_XBOOTH/XSEL02/B_XBOOTH/Xsel02/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa27/Xyb1/M10 N_XADDER/XA27/XYB1/N004_XADDER/Xa27/Xyb1/M10_d
+ N_XADDER/PP7_XADDER/Xa27/Xyb1/M10_g N_GND_XADDER/Xa27/Xyb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=9.24e-14 AS=2.244e-13
+ PD=4.2e-07 PS=1.46e-06
mXCSA/Xdffa3/M9 N_XCSA/XDFFA3/P003_XCSA/Xdffa3/M9_d
+ N_XCSA/XDFFA3/N1_XCSA/Xdffa3/M9_g N_GND_XCSA/Xdffa3/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/Xdffa16/M9 N_XCSA/XDFFA16/P003_XCSA/Xdffa16/M9_d
+ N_XCSA/XDFFA16/N1_XCSA/Xdffa16/M9_g N_GND_XCSA/Xdffa16/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mX02/xd27/M11 N_OUT[6]_X02/xd27/M11_d N_X02/XD27/N3_X02/xd27/M11_g
+ N_GND_X02/xd27/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/X_LV3_FA2/M25 N_XCSA/LV3_S[4]_XCSA/X_LV3_FA2/M25_d
+ N_XCSA/X_LV3_FA2/_SUM_XCSA/X_LV3_FA2/M25_g N_GND_XCSA/X_LV3_FA2/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xdffb2/M11 N_XBOOTH/B_D[2]_XBOOTH/Xdffb2/M11_d
+ N_XBOOTH/XDFFB2/N3_XBOOTH/Xdffb2/M11_g N_GND_XBOOTH/Xdffb2/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXADDER/Xa37/Xao2/M37 N_XADDER/XA37/XAO2/N008_XADDER/Xa37/Xao2/M37_d
+ N_XADDER/XA37/OUT1_XADDER/Xa37/Xao2/M37_g N_GND_XADDER/Xa37/Xao2/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel22/M11 N_XBOOTH/XSEL22/N004_XBOOTH/Xsel22/M11_d
+ N_XBOOTH/XSEL22/B_XBOOTH/Xsel22/M11_g N_A_D[5]_XBOOTH/Xsel22/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel12/M11 N_XBOOTH/XSEL12/N004_XBOOTH/Xsel12/M11_d
+ N_XBOOTH/XSEL12/B_XBOOTH/Xsel12/M11_g N_A_D[3]_XBOOTH/Xsel12/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel02/M11 N_XBOOTH/XSEL02/N004_XBOOTH/Xsel02/M11_d
+ N_XBOOTH/XSEL02/B_XBOOTH/Xsel02/M11_g N_A_D[1]_XBOOTH/Xsel02/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/Xdffa3/M11 N_C[4]_XCSA/Xdffa3/M11_d N_XCSA/XDFFA3/N3_XCSA/Xdffa3/M11_g
+ N_GND_XCSA/Xdffa3/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/Xdffa16/M11 N_S[4]_XCSA/Xdffa16/M11_d N_XCSA/XDFFA16/N3_XCSA/Xdffa16/M11_g
+ N_GND_XCSA/Xdffa16/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXADDER/Xa06/Xrb1/Xand1/M16 N_XADDER/G5_XADDER/Xa06/Xrb1/Xand1/M16_d
+ N_XADDER/XA06/XRB1/N003_XADDER/Xa06/Xrb1/Xand1/M16_g
+ N_GND_XADDER/Xa06/Xrb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA4/X_xor/M2 N_XCSA/X_LV2_HA4/X_XOR/N002_XCSA/X_LV2_HA4/X_xor/M2_d
+ N_XCSA/LV1_C[6]_XCSA/X_LV2_HA4/X_xor/M2_g
+ N_XCSA/LV1_S[6]_XCSA/X_LV2_HA4/X_xor/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13 PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA4/M11 N_XCSA/X_LV2_HA4/P001_XCSA/X_LV2_HA4/M11_d
+ N_XCSA/LV1_C[6]_XCSA/X_LV2_HA4/M11_g N_GND_XCSA/X_LV2_HA4/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV1_FA2/M19 N_XCSA/X_LV1_FA2/N004_XCSA/X_LV1_FA2/M19_d
+ N_PP0[6]_XCSA/X_LV1_FA2/M19_g N_GND_XCSA/X_LV1_FA2/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA2/M24 N_XCSA/X_LV1_FA2/P006_XCSA/X_LV1_FA2/M24_d
+ N_PP0[6]_XCSA/X_LV1_FA2/M24_g N_GND_XCSA/X_LV1_FA2/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA2/M14 N_XCSA/X_LV1_FA2/P004_XCSA/X_LV1_FA2/M14_d
+ N_PP0[6]_XCSA/X_LV1_FA2/M14_g N_GND_XCSA/X_LV1_FA2/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA2/M16 N_XCSA/X_LV1_FA2/N003_XCSA/X_LV1_FA2/M16_d
+ N_PP0[6]_XCSA/X_LV1_FA2/M16_g N_GND_XCSA/X_LV1_FA2/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA2/M26 N_XCSA/LV3_C[5]_XCSA/X_LV3_FA2/M26_d
+ N_XCSA/X_LV3_FA2/_COUT_XCSA/X_LV3_FA2/M26_g N_GND_XCSA/X_LV3_FA2/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa37/Xao2/M38 N_XADDER/XA37/XAO2/N008_XADDER/Xa37/Xao2/M38_d
+ N_XADDER/GGG7_XADDER/Xa37/Xao2/M38_g N_GND_XADDER/Xa37/Xao2/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa27/Xyb2/M10 N_XADDER/XA27/XYB2/N004_XADDER/Xa27/Xyb2/M10_d
+ N_XADDER/PP7_XADDER/Xa27/Xyb2/M10_g N_GND_XADDER/Xa27/Xyb2/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXBOOTH/Xsel22/M13 N_PP2[2]_XBOOTH/Xsel22/M13_d
+ N_XBOOTH/XSEL22/N004_XBOOTH/Xsel22/M13_g N_GND_XBOOTH/Xsel22/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel12/M13 N_PP1[2]_XBOOTH/Xsel12/M13_d
+ N_XBOOTH/XSEL12/N004_XBOOTH/Xsel12/M13_g N_GND_XBOOTH/Xsel12/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel02/M13 N_PP0[2]_XBOOTH/Xsel02/M13_d
+ N_XBOOTH/XSEL02/N004_XBOOTH/Xsel02/M13_g N_GND_XBOOTH/Xsel02/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA2/M21 N_XCSA/X_LV3_FA2/_SUM_XCSA/X_LV3_FA2/M21_d
+ N_XCSA/X_LV3_FA2/_COUT_XCSA/X_LV3_FA2/M21_g
+ N_XCSA/X_LV3_FA2/N004_XCSA/X_LV3_FA2/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXCSA/X_LV2_HA4/X_xor/M1 N_XCSA/X_LV2_HA4/X_XOR/N002_XCSA/X_LV2_HA4/X_xor/M1_d
+ N_XCSA/LV1_S[6]_XCSA/X_LV2_HA4/X_xor/M1_g
+ N_XCSA/LV1_C[6]_XCSA/X_LV2_HA4/X_xor/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_HA4/M12 N_XCSA/X_LV2_HA4/N001_XCSA/X_LV2_HA4/M12_d
+ N_XCSA/LV1_S[6]_XCSA/X_LV2_HA4/M12_g
+ N_XCSA/X_LV2_HA4/P001_XCSA/X_LV2_HA4/M12_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA2/M20 N_XCSA/X_LV1_FA2/N004_XCSA/X_LV1_FA2/M20_d
+ N_PP1[4]_XCSA/X_LV1_FA2/M20_g N_GND_XCSA/X_LV1_FA2/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV1_FA2/M23 N_XCSA/X_LV1_FA2/P005_XCSA/X_LV1_FA2/M23_d
+ N_PP1[4]_XCSA/X_LV1_FA2/M23_g N_XCSA/X_LV1_FA2/P006_XCSA/X_LV1_FA2/M23_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA2/M13 N_XCSA/X_LV1_FA2/_COUT_XCSA/X_LV1_FA2/M13_d
+ N_PP1[4]_XCSA/X_LV1_FA2/M13_g N_XCSA/X_LV1_FA2/P004_XCSA/X_LV1_FA2/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA2/M17 N_XCSA/X_LV1_FA2/N003_XCSA/X_LV1_FA2/M17_d
+ N_PP1[4]_XCSA/X_LV1_FA2/M17_g N_GND_XCSA/X_LV1_FA2/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXADDER/Xa27/Xyb2/M9 N_XADDER/XA27/XYB2/N003_XADDER/Xa27/Xyb2/M9_d
+ N_XADDER/GG5_XADDER/Xa27/Xyb2/M9_g
+ N_XADDER/XA27/XYB2/N004_XADDER/Xa27/Xyb2/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=6.16e-14 PD=1.74e-06 PS=2.8e-07
mXCSA/Xdffa4/M3 N_XCSA/XDFFA4/N0_XCSA/Xdffa4/M3_d
+ N_XCSA/LV3_C[5]_XCSA/Xdffa4/M3_g N_GND_XCSA/Xdffa4/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa17/M3 N_XCSA/XDFFA17/N0_XCSA/Xdffa17/M3_d
+ N_XCSA/LV3_S[5]_XCSA/Xdffa17/M3_g N_GND_XCSA/Xdffa17/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA2/M18 N_XCSA/X_LV1_FA2/N004_XCSA/X_LV1_FA2/M18_d
+ N_PP2[2]_XCSA/X_LV1_FA2/M18_g N_GND_XCSA/X_LV1_FA2/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV1_FA2/M22 N_XCSA/X_LV1_FA2/_SUM_XCSA/X_LV1_FA2/M22_d
+ N_PP2[2]_XCSA/X_LV1_FA2/M22_g N_XCSA/X_LV1_FA2/P005_XCSA/X_LV1_FA2/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV1_FA2/M15 N_XCSA/X_LV1_FA2/_COUT_XCSA/X_LV1_FA2/M15_d
+ N_PP2[2]_XCSA/X_LV1_FA2/M15_g N_XCSA/X_LV1_FA2/N003_XCSA/X_LV1_FA2/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV3_FA2/M18 N_XCSA/X_LV3_FA2/N004_XCSA/X_LV3_FA2/M18_d
+ N_CACC[4]_XCSA/X_LV3_FA2/M18_g N_GND_XCSA/X_LV3_FA2/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA2/M22 N_XCSA/X_LV3_FA2/_SUM_XCSA/X_LV3_FA2/M22_d
+ N_CACC[4]_XCSA/X_LV3_FA2/M22_g N_XCSA/X_LV3_FA2/P005_XCSA/X_LV3_FA2/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV3_FA2/M15 N_XCSA/X_LV3_FA2/_COUT_XCSA/X_LV3_FA2/M15_d
+ N_CACC[4]_XCSA/X_LV3_FA2/M15_g N_XCSA/X_LV3_FA2/N003_XCSA/X_LV3_FA2/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXADDER/Xa37/Xao2/Xor1/M16 N_XADDER/GOUT7_XADDER/Xa37/Xao2/Xor1/M16_d
+ N_XADDER/XA37/XAO2/N008_XADDER/Xa37/Xao2/Xor1/M16_g
+ N_GND_XADDER/Xa37/Xao2/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa17/Xyb1/Xand1/M16 N_XADDER/PP7_XADDER/Xa17/Xyb1/Xand1/M16_d
+ N_XADDER/XA17/XYB1/N003_XADDER/Xa17/Xyb1/Xand1/M16_g
+ N_GND_XADDER/Xa17/Xyb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa07/Xrb2/M3 N_XADDER/P6_XADDER/Xa07/Xrb2/M3_d
+ N_XADDER/XA07/XRB2/N002_XADDER/Xa07/Xrb2/M3_g N_GND_XADDER/Xa07/Xrb2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa4/M6 N_XCSA/XDFFA4/P002_XCSA/Xdffa4/M6_d N_CLK_XCSA/Xdffa4/M6_g
+ N_GND_XCSA/Xdffa4/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/Xdffa17/M6 N_XCSA/XDFFA17/P002_XCSA/Xdffa17/M6_d N_CLK_XCSA/Xdffa17/M6_g
+ N_GND_XCSA/Xdffa17/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/X_LV2_HA4/X_xor/M3 N_XCSA/LV2_S[6]_XCSA/X_LV2_HA4/X_xor/M3_d
+ N_XCSA/X_LV2_HA4/X_XOR/N002_XCSA/X_LV2_HA4/X_xor/M3_g
+ N_GND_XCSA/X_LV2_HA4/X_xor/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA4/M14 N_XCSA/LV2_C[7]_XCSA/X_LV2_HA4/M14_d
+ N_XCSA/X_LV2_HA4/N001_XCSA/X_LV2_HA4/M14_g N_GND_XCSA/X_LV2_HA4/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA2/M20 N_XCSA/X_LV3_FA2/N004_XCSA/X_LV3_FA2/M20_d
+ N_XCSA/LV2_S[4]_XCSA/X_LV3_FA2/M20_g N_GND_XCSA/X_LV3_FA2/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA2/M23 N_XCSA/X_LV3_FA2/P005_XCSA/X_LV3_FA2/M23_d
+ N_XCSA/LV2_S[4]_XCSA/X_LV3_FA2/M23_g
+ N_XCSA/X_LV3_FA2/P006_XCSA/X_LV3_FA2/M23_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA2/M13 N_XCSA/X_LV3_FA2/_COUT_XCSA/X_LV3_FA2/M13_d
+ N_XCSA/LV2_S[4]_XCSA/X_LV3_FA2/M13_g
+ N_XCSA/X_LV3_FA2/P004_XCSA/X_LV3_FA2/M13_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA2/M17 N_XCSA/X_LV3_FA2/N003_XCSA/X_LV3_FA2/M17_d
+ N_XCSA/LV2_S[4]_XCSA/X_LV3_FA2/M17_g N_GND_XCSA/X_LV3_FA2/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA2/M21 N_XCSA/X_LV1_FA2/_SUM_XCSA/X_LV1_FA2/M21_d
+ N_XCSA/X_LV1_FA2/_COUT_XCSA/X_LV1_FA2/M21_g
+ N_XCSA/X_LV1_FA2/N004_XCSA/X_LV1_FA2/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXADDER/Xa27/Xyb2/Xand1/M16 N_XADDER/XA27/T1_XADDER/Xa27/Xyb2/Xand1/M16_d
+ N_XADDER/XA27/XYB2/N003_XADDER/Xa27/Xyb2/Xand1/M16_g
+ N_GND_XADDER/Xa27/Xyb2/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa4/M5 N_XCSA/XDFFA4/N1_XCSA/Xdffa4/M5_d
+ N_XCSA/XDFFA4/N0_XCSA/Xdffa4/M5_g N_XCSA/XDFFA4/P002_XCSA/Xdffa4/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa17/M5 N_XCSA/XDFFA17/N1_XCSA/Xdffa17/M5_d
+ N_XCSA/XDFFA17/N0_XCSA/Xdffa17/M5_g N_XCSA/XDFFA17/P002_XCSA/Xdffa17/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel23/M2 N_noxref_2198_XBOOTH/Xsel23/M2_d
+ N_XBOOTH/B_D[2]_XBOOTH/Xsel23/M2_g N_GND_XBOOTH/Xsel23/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel13/M2 N_noxref_2199_XBOOTH/Xsel13/M2_d
+ N_XBOOTH/B_D[2]_XBOOTH/Xsel13/M2_g N_GND_XBOOTH/Xsel13/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel03/M2 N_noxref_2200_XBOOTH/Xsel03/M2_d
+ N_XBOOTH/B_D[2]_XBOOTH/Xsel03/M2_g N_GND_XBOOTH/Xsel03/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA2/M26 N_XCSA/LV1_C[7]_XCSA/X_LV1_FA2/M26_d
+ N_XCSA/X_LV1_FA2/_COUT_XCSA/X_LV1_FA2/M26_g N_GND_XCSA/X_LV1_FA2/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA2/M19 N_XCSA/X_LV3_FA2/N004_XCSA/X_LV3_FA2/M19_d
+ N_XCSA/LV2_C[4]_XCSA/X_LV3_FA2/M19_g N_GND_XCSA/X_LV3_FA2/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA2/M24 N_XCSA/X_LV3_FA2/P006_XCSA/X_LV3_FA2/M24_d
+ N_XCSA/LV2_C[4]_XCSA/X_LV3_FA2/M24_g N_GND_XCSA/X_LV3_FA2/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA2/M14 N_XCSA/X_LV3_FA2/P004_XCSA/X_LV3_FA2/M14_d
+ N_XCSA/LV2_C[4]_XCSA/X_LV3_FA2/M14_g N_GND_XCSA/X_LV3_FA2/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA2/M16 N_XCSA/X_LV3_FA2/N003_XCSA/X_LV3_FA2/M16_d
+ N_XCSA/LV2_C[4]_XCSA/X_LV3_FA2/M16_g N_GND_XCSA/X_LV3_FA2/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa17/Xyb1/M9 N_XADDER/XA17/XYB1/N003_XADDER/Xa17/Xyb1/M9_d
+ N_XADDER/P6_XADDER/Xa17/Xyb1/M9_g
+ N_XADDER/XA17/XYB1/N004_XADDER/Xa17/Xyb1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=9.24e-14 PD=1.44e-06 PS=4.2e-07
mXADDER/Xa07/Xrb2/M1 N_XADDER/XA07/XRB2/N002_XADDER/Xa07/Xrb2/M1_d
+ N_C[6]_XADDER/Xa07/Xrb2/M1_g N_S[6]_XADDER/Xa07/Xrb2/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel23/M1 N_XBOOTH/XSEL23/N002_XBOOTH/Xsel23/M1_d
+ N_XBOOTH/D2_XBOOTH/Xsel23/M1_g N_noxref_2198_XBOOTH/Xsel23/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel13/M1 N_XBOOTH/XSEL13/N002_XBOOTH/Xsel13/M1_d
+ N_XBOOTH/D1_XBOOTH/Xsel13/M1_g N_noxref_2199_XBOOTH/Xsel13/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel03/M1 N_XBOOTH/XSEL03/N002_XBOOTH/Xsel03/M1_d
+ N_XBOOTH/D0_XBOOTH/Xsel03/M1_g N_noxref_2200_XBOOTH/Xsel03/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXADDER/Xa17/Xyb1/M10 N_XADDER/XA17/XYB1/N004_XADDER/Xa17/Xyb1/M10_d
+ N_XADDER/P7_XADDER/Xa17/Xyb1/M10_g N_GND_XADDER/Xa17/Xyb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=9.24e-14 AS=2.244e-13
+ PD=4.2e-07 PS=1.46e-06
mXCSA/X_LV1_FA2/M25 N_XCSA/LV1_S[6]_XCSA/X_LV1_FA2/M25_d
+ N_XCSA/X_LV1_FA2/_SUM_XCSA/X_LV1_FA2/M25_g N_GND_XCSA/X_LV1_FA2/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xdffb3/M3 N_XBOOTH/XDFFB3/N0_XBOOTH/Xdffb3/M3_d
+ N_B[3]_XBOOTH/Xdffb3/M3_g N_GND_XBOOTH/Xdffb3/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa07/Xrb2/M2 N_XADDER/XA07/XRB2/N002_XADDER/Xa07/Xrb2/M2_d
+ N_S[6]_XADDER/Xa07/Xrb2/M2_g N_C[6]_XADDER/Xa07/Xrb2/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXADDER/Xa27/Xyb3/M37 N_XADDER/XA27/XYB3/N008_XADDER/Xa27/Xyb3/M37_d
+ N_XADDER/XA27/T1_XADDER/Xa27/Xyb3/M37_g N_GND_XADDER/Xa27/Xyb3/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa4/M8 N_XCSA/XDFFA4/N3_XCSA/Xdffa4/M8_d N_CLK_XCSA/Xdffa4/M8_g
+ N_XCSA/XDFFA4/P003_XCSA/Xdffa4/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa17/M8 N_XCSA/XDFFA17/N3_XCSA/Xdffa17/M8_d N_CLK_XCSA/Xdffa17/M8_g
+ N_XCSA/XDFFA17/P003_XCSA/Xdffa17/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel23/M3 N_XBOOTH/XSEL23/N002_XBOOTH/Xsel23/M3_d
+ N_XBOOTH/S2_XBOOTH/Xsel23/M3_g N_noxref_2204_XBOOTH/Xsel23/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel13/M3 N_XBOOTH/XSEL13/N002_XBOOTH/Xsel13/M3_d
+ N_XBOOTH/S1_XBOOTH/Xsel13/M3_g N_noxref_2205_XBOOTH/Xsel13/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel03/M3 N_XBOOTH/XSEL03/N002_XBOOTH/Xsel03/M3_d
+ N_XBOOTH/S0_XBOOTH/Xsel03/M3_g N_noxref_2206_XBOOTH/Xsel03/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXCSA/Xdffa4/M9 N_XCSA/XDFFA4/P003_XCSA/Xdffa4/M9_d
+ N_XCSA/XDFFA4/N1_XCSA/Xdffa4/M9_g N_GND_XCSA/Xdffa4/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/Xdffa17/M9 N_XCSA/XDFFA17/P003_XCSA/Xdffa17/M9_d
+ N_XCSA/XDFFA17/N1_XCSA/Xdffa17/M9_g N_GND_XCSA/Xdffa17/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/X_LV3_FA3/M25 N_XCSA/LV3_S[5]_XCSA/X_LV3_FA3/M25_d
+ N_XCSA/X_LV3_FA3/_SUM_XCSA/X_LV3_FA3/M25_g N_GND_XCSA/X_LV3_FA3/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xdffb3/M6 N_XBOOTH/XDFFB3/P002_XBOOTH/Xdffb3/M6_d
+ N_CLK_XBOOTH/Xdffb3/M6_g N_GND_XBOOTH/Xdffb3/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXADDER/Xa27/Xyb3/M38 N_XADDER/XA27/XYB3/N008_XADDER/Xa27/Xyb3/M38_d
+ N_XADDER/GG7_XADDER/Xa27/Xyb3/M38_g N_GND_XADDER/Xa27/Xyb3/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel23/M4 N_noxref_2204_XBOOTH/Xsel23/M4_d
+ N_XBOOTH/B_D[3]_XBOOTH/Xsel23/M4_g N_GND_XBOOTH/Xsel23/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel13/M4 N_noxref_2205_XBOOTH/Xsel13/M4_d
+ N_XBOOTH/B_D[3]_XBOOTH/Xsel13/M4_g N_GND_XBOOTH/Xsel13/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel03/M4 N_noxref_2206_XBOOTH/Xsel03/M4_d
+ N_XBOOTH/B_D[3]_XBOOTH/Xsel03/M4_g N_GND_XBOOTH/Xsel03/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xdffb3/M5 N_XBOOTH/XDFFB3/N1_XBOOTH/Xdffb3/M5_d
+ N_XBOOTH/XDFFB3/N0_XBOOTH/Xdffb3/M5_g N_XBOOTH/XDFFB3/P002_XBOOTH/Xdffb3/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa17/Xyb2/M10 N_XADDER/XA17/XYB2/N004_XADDER/Xa17/Xyb2/M10_d
+ N_XADDER/P7_XADDER/Xa17/Xyb2/M10_g N_GND_XADDER/Xa17/Xyb2/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXCSA/X_LV3_FA3/M26 N_XCSA/LV3_C[6]_XCSA/X_LV3_FA3/M26_d
+ N_XCSA/X_LV3_FA3/_COUT_XCSA/X_LV3_FA3/M26_g N_GND_XCSA/X_LV3_FA3/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa07/Xrb1/M10 N_XADDER/XA07/XRB1/N004_XADDER/Xa07/Xrb1/M10_d
+ N_S[6]_XADDER/Xa07/Xrb1/M10_g N_GND_XADDER/Xa07/Xrb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXCSA/Xdffa4/M11 N_C[5]_XCSA/Xdffa4/M11_d N_XCSA/XDFFA4/N3_XCSA/Xdffa4/M11_g
+ N_GND_XCSA/Xdffa4/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/Xdffa17/M11 N_S[5]_XCSA/Xdffa17/M11_d N_XCSA/XDFFA17/N3_XCSA/Xdffa17/M11_g
+ N_GND_XCSA/Xdffa17/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXBOOTH/Xsel23/M5 N_XBOOTH/XSEL23/B_XBOOTH/Xsel23/M5_d
+ N_XBOOTH/XSEL23/N002_XBOOTH/Xsel23/M5_g N_GND_XBOOTH/Xsel23/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel13/M5 N_XBOOTH/XSEL13/B_XBOOTH/Xsel13/M5_d
+ N_XBOOTH/XSEL13/N002_XBOOTH/Xsel13/M5_g N_GND_XBOOTH/Xsel13/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel03/M5 N_XBOOTH/XSEL03/B_XBOOTH/Xsel03/M5_d
+ N_XBOOTH/XSEL03/N002_XBOOTH/Xsel03/M5_g N_GND_XBOOTH/Xsel03/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa17/Xyb2/M9 N_XADDER/XA17/XYB2/N003_XADDER/Xa17/Xyb2/M9_d
+ N_XADDER/G6_XADDER/Xa17/Xyb2/M9_g
+ N_XADDER/XA17/XYB2/N004_XADDER/Xa17/Xyb2/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=6.16e-14 PD=1.74e-06 PS=2.8e-07
mXADDER/Xa07/Xrb1/M9 N_XADDER/XA07/XRB1/N003_XADDER/Xa07/Xrb1/M9_d
+ N_C[6]_XADDER/Xa07/Xrb1/M9_g N_XADDER/XA07/XRB1/N004_XADDER/Xa07/Xrb1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14
+ PD=1.44e-06 PS=2.8e-07
mXCSA/X_LV3_FA3/M21 N_XCSA/X_LV3_FA3/_SUM_XCSA/X_LV3_FA3/M21_d
+ N_XCSA/X_LV3_FA3/_COUT_XCSA/X_LV3_FA3/M21_g
+ N_XCSA/X_LV3_FA3/N004_XCSA/X_LV3_FA3/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXCSA/X_LV1_FA3/M19 N_XCSA/X_LV1_FA3/N004_XCSA/X_LV1_FA3/M19_d
+ N_PP0[6]_XCSA/X_LV1_FA3/M19_g N_GND_XCSA/X_LV1_FA3/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA3/M24 N_XCSA/X_LV1_FA3/P006_XCSA/X_LV1_FA3/M24_d
+ N_PP0[6]_XCSA/X_LV1_FA3/M24_g N_GND_XCSA/X_LV1_FA3/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA3/M14 N_XCSA/X_LV1_FA3/P004_XCSA/X_LV1_FA3/M14_d
+ N_PP0[6]_XCSA/X_LV1_FA3/M14_g N_GND_XCSA/X_LV1_FA3/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA3/M16 N_XCSA/X_LV1_FA3/N003_XCSA/X_LV1_FA3/M16_d
+ N_PP0[6]_XCSA/X_LV1_FA3/M16_g N_GND_XCSA/X_LV1_FA3/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa27/Xyb3/Xor1/M16 N_XADDER/GGG7_XADDER/Xa27/Xyb3/Xor1/M16_d
+ N_XADDER/XA27/XYB3/N008_XADDER/Xa27/Xyb3/Xor1/M16_g
+ N_GND_XADDER/Xa27/Xyb3/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa76/M3 N_OUT1[6]_XADDER/Xa76/M3_d N_XADDER/XA76/N002_XADDER/Xa76/M3_g
+ N_GND_XADDER/Xa76/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd29/M3 N_X02/XD29/N0_X02/xd29/M3_d N_OUT1[8]_X02/xd29/M3_g
+ N_GND_X02/xd29/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xdffb3/M8 N_XBOOTH/XDFFB3/N3_XBOOTH/Xdffb3/M8_d N_CLK_XBOOTH/Xdffb3/M8_g
+ N_XBOOTH/XDFFB3/P003_XBOOTH/Xdffb3/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV2_HA5/X_xor/M2 N_XCSA/X_LV2_HA5/X_XOR/N002_XCSA/X_LV2_HA5/X_xor/M2_d
+ N_XCSA/LV1_C[7]_XCSA/X_LV2_HA5/X_xor/M2_g
+ N_XCSA/LV1_S[7]_XCSA/X_LV2_HA5/X_xor/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13 PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA5/M11 N_XCSA/X_LV2_HA5/P001_XCSA/X_LV2_HA5/M11_d
+ N_XCSA/LV1_C[7]_XCSA/X_LV2_HA5/M11_g N_GND_XCSA/X_LV2_HA5/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV1_FA3/M20 N_XCSA/X_LV1_FA3/N004_XCSA/X_LV1_FA3/M20_d
+ N_PP1[5]_XCSA/X_LV1_FA3/M20_g N_GND_XCSA/X_LV1_FA3/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV1_FA3/M23 N_XCSA/X_LV1_FA3/P005_XCSA/X_LV1_FA3/M23_d
+ N_PP1[5]_XCSA/X_LV1_FA3/M23_g N_XCSA/X_LV1_FA3/P006_XCSA/X_LV1_FA3/M23_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA3/M13 N_XCSA/X_LV1_FA3/_COUT_XCSA/X_LV1_FA3/M13_d
+ N_PP1[5]_XCSA/X_LV1_FA3/M13_g N_XCSA/X_LV1_FA3/P004_XCSA/X_LV1_FA3/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA3/M17 N_XCSA/X_LV1_FA3/N003_XCSA/X_LV1_FA3/M17_d
+ N_PP1[5]_XCSA/X_LV1_FA3/M17_g N_GND_XCSA/X_LV1_FA3/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA3/M18 N_XCSA/X_LV3_FA3/N004_XCSA/X_LV3_FA3/M18_d
+ N_CACC[5]_XCSA/X_LV3_FA3/M18_g N_GND_XCSA/X_LV3_FA3/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA3/M22 N_XCSA/X_LV3_FA3/_SUM_XCSA/X_LV3_FA3/M22_d
+ N_CACC[5]_XCSA/X_LV3_FA3/M22_g N_XCSA/X_LV3_FA3/P005_XCSA/X_LV3_FA3/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV3_FA3/M15 N_XCSA/X_LV3_FA3/_COUT_XCSA/X_LV3_FA3/M15_d
+ N_CACC[5]_XCSA/X_LV3_FA3/M15_g N_XCSA/X_LV3_FA3/N003_XCSA/X_LV3_FA3/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXBOOTH/Xdffb3/M9 N_XBOOTH/XDFFB3/P003_XBOOTH/Xdffb3/M9_d
+ N_XBOOTH/XDFFB3/N1_XBOOTH/Xdffb3/M9_g N_GND_XBOOTH/Xdffb3/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/Xdffa5/M3 N_XCSA/XDFFA5/N0_XCSA/Xdffa5/M3_d
+ N_XCSA/LV3_C[6]_XCSA/Xdffa5/M3_g N_GND_XCSA/Xdffa5/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa18/M3 N_XCSA/XDFFA18/N0_XCSA/Xdffa18/M3_d
+ N_XCSA/LV3_S[6]_XCSA/Xdffa18/M3_g N_GND_XCSA/Xdffa18/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd29/M6 N_X02/XD29/P002_X02/xd29/M6_d N_CLK_X02/xd29/M6_g
+ N_GND_X02/xd29/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/X_LV2_HA5/X_xor/M1 N_XCSA/X_LV2_HA5/X_XOR/N002_XCSA/X_LV2_HA5/X_xor/M1_d
+ N_XCSA/LV1_S[7]_XCSA/X_LV2_HA5/X_xor/M1_g
+ N_XCSA/LV1_C[7]_XCSA/X_LV2_HA5/X_xor/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_HA5/M12 N_XCSA/X_LV2_HA5/N001_XCSA/X_LV2_HA5/M12_d
+ N_XCSA/LV1_S[7]_XCSA/X_LV2_HA5/M12_g
+ N_XCSA/X_LV2_HA5/P001_XCSA/X_LV2_HA5/M12_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXADDER/Xa17/Xyb2/Xand1/M16 N_XADDER/XA17/T1_XADDER/Xa17/Xyb2/Xand1/M16_d
+ N_XADDER/XA17/XYB2/N003_XADDER/Xa17/Xyb2/Xand1/M16_g
+ N_GND_XADDER/Xa17/Xyb2/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa07/Xrb1/Xand1/M16 N_XADDER/G6_XADDER/Xa07/Xrb1/Xand1/M16_d
+ N_XADDER/XA07/XRB1/N003_XADDER/Xa07/Xrb1/Xand1/M16_g
+ N_GND_XADDER/Xa07/Xrb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd29/M5 N_X02/XD29/N1_X02/xd29/M5_d N_X02/XD29/N0_X02/xd29/M5_g
+ N_X02/XD29/P002_X02/xd29/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV1_FA3/M18 N_XCSA/X_LV1_FA3/N004_XCSA/X_LV1_FA3/M18_d
+ N_PP2[3]_XCSA/X_LV1_FA3/M18_g N_GND_XCSA/X_LV1_FA3/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV1_FA3/M22 N_XCSA/X_LV1_FA3/_SUM_XCSA/X_LV1_FA3/M22_d
+ N_PP2[3]_XCSA/X_LV1_FA3/M22_g N_XCSA/X_LV1_FA3/P005_XCSA/X_LV1_FA3/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV1_FA3/M15 N_XCSA/X_LV1_FA3/_COUT_XCSA/X_LV1_FA3/M15_d
+ N_PP2[3]_XCSA/X_LV1_FA3/M15_g N_XCSA/X_LV1_FA3/N003_XCSA/X_LV1_FA3/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV3_FA3/M20 N_XCSA/X_LV3_FA3/N004_XCSA/X_LV3_FA3/M20_d
+ N_XCSA/LV2_S[5]_XCSA/X_LV3_FA3/M20_g N_GND_XCSA/X_LV3_FA3/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA3/M23 N_XCSA/X_LV3_FA3/P005_XCSA/X_LV3_FA3/M23_d
+ N_XCSA/LV2_S[5]_XCSA/X_LV3_FA3/M23_g
+ N_XCSA/X_LV3_FA3/P006_XCSA/X_LV3_FA3/M23_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA3/M13 N_XCSA/X_LV3_FA3/_COUT_XCSA/X_LV3_FA3/M13_d
+ N_XCSA/LV2_S[5]_XCSA/X_LV3_FA3/M13_g
+ N_XCSA/X_LV3_FA3/P004_XCSA/X_LV3_FA3/M13_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA3/M17 N_XCSA/X_LV3_FA3/N003_XCSA/X_LV3_FA3/M17_d
+ N_XCSA/LV2_S[5]_XCSA/X_LV3_FA3/M17_g N_GND_XCSA/X_LV3_FA3/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXBOOTH/Xsel23/M12 N_XBOOTH/XSEL23/N004_XBOOTH/Xsel23/M12_d
+ N_A_D[5]_XBOOTH/Xsel23/M12_g N_XBOOTH/XSEL23/B_XBOOTH/Xsel23/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel13/M12 N_XBOOTH/XSEL13/N004_XBOOTH/Xsel13/M12_d
+ N_A_D[3]_XBOOTH/Xsel13/M12_g N_XBOOTH/XSEL13/B_XBOOTH/Xsel13/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel03/M12 N_XBOOTH/XSEL03/N004_XBOOTH/Xsel03/M12_d
+ N_A_D[1]_XBOOTH/Xsel03/M12_g N_XBOOTH/XSEL03/B_XBOOTH/Xsel03/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/Xdffa5/M6 N_XCSA/XDFFA5/P002_XCSA/Xdffa5/M6_d N_CLK_XCSA/Xdffa5/M6_g
+ N_GND_XCSA/Xdffa5/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/Xdffa18/M6 N_XCSA/XDFFA18/P002_XCSA/Xdffa18/M6_d N_CLK_XCSA/Xdffa18/M6_g
+ N_GND_XCSA/Xdffa18/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXADDER/Xa66/Xao1/M9 N_XADDER/XA66/XAO1/N003_XADDER/Xa66/Xao1/M9_d
+ N_XADDER/GX5[0]_XADDER/Xa66/Xao1/M9_g
+ N_XADDER/XA66/XAO1/N004_XADDER/Xa66/Xao1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14 PD=1.44e-06 PS=2.8e-07
mXBOOTH/Xdffb3/M11 N_XBOOTH/B_D[3]_XBOOTH/Xdffb3/M11_d
+ N_XBOOTH/XDFFB3/N3_XBOOTH/Xdffb3/M11_g N_GND_XBOOTH/Xdffb3/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXCSA/Xdffa5/M5 N_XCSA/XDFFA5/N1_XCSA/Xdffa5/M5_d
+ N_XCSA/XDFFA5/N0_XCSA/Xdffa5/M5_g N_XCSA/XDFFA5/P002_XCSA/Xdffa5/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa18/M5 N_XCSA/XDFFA18/N1_XCSA/Xdffa18/M5_d
+ N_XCSA/XDFFA18/N0_XCSA/Xdffa18/M5_g N_XCSA/XDFFA18/P002_XCSA/Xdffa18/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa76/M1 N_XADDER/XA76/N002_XADDER/Xa76/M1_d N_XADDER/P6_XADDER/Xa76/M1_g
+ N_XADDER/GX5[0]_XADDER/Xa76/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=2.332e-13 PD=5.4e-07 PS=1.5e-06
mXADDER/Xa66/Xao1/M10 N_XADDER/XA66/XAO1/N004_XADDER/Xa66/Xao1/M10_d
+ N_XADDER/P6_XADDER/Xa66/Xao1/M10_g N_GND_XADDER/Xa66/Xao1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.86e-13
+ PD=2.8e-07 PS=1.74e-06
mXCSA/X_LV3_FA3/M19 N_XCSA/X_LV3_FA3/N004_XCSA/X_LV3_FA3/M19_d
+ N_XCSA/LV2_C[5]_XCSA/X_LV3_FA3/M19_g N_GND_XCSA/X_LV3_FA3/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA3/M24 N_XCSA/X_LV3_FA3/P006_XCSA/X_LV3_FA3/M24_d
+ N_XCSA/LV2_C[5]_XCSA/X_LV3_FA3/M24_g N_GND_XCSA/X_LV3_FA3/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA3/M14 N_XCSA/X_LV3_FA3/P004_XCSA/X_LV3_FA3/M14_d
+ N_XCSA/LV2_C[5]_XCSA/X_LV3_FA3/M14_g N_GND_XCSA/X_LV3_FA3/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA3/M16 N_XCSA/X_LV3_FA3/N003_XCSA/X_LV3_FA3/M16_d
+ N_XCSA/LV2_C[5]_XCSA/X_LV3_FA3/M16_g N_GND_XCSA/X_LV3_FA3/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA3/M21 N_XCSA/X_LV1_FA3/_SUM_XCSA/X_LV1_FA3/M21_d
+ N_XCSA/X_LV1_FA3/_COUT_XCSA/X_LV1_FA3/M21_g
+ N_XCSA/X_LV1_FA3/N004_XCSA/X_LV1_FA3/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXBOOTH/Xsel23/M11 N_XBOOTH/XSEL23/N004_XBOOTH/Xsel23/M11_d
+ N_XBOOTH/XSEL23/B_XBOOTH/Xsel23/M11_g N_A_D[5]_XBOOTH/Xsel23/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel13/M11 N_XBOOTH/XSEL13/N004_XBOOTH/Xsel13/M11_d
+ N_XBOOTH/XSEL13/B_XBOOTH/Xsel13/M11_g N_A_D[3]_XBOOTH/Xsel13/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel03/M11 N_XBOOTH/XSEL03/N004_XBOOTH/Xsel03/M11_d
+ N_XBOOTH/XSEL03/B_XBOOTH/Xsel03/M11_g N_A_D[1]_XBOOTH/Xsel03/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_HA5/X_xor/M3 N_XCSA/LV2_S[7]_XCSA/X_LV2_HA5/X_xor/M3_d
+ N_XCSA/X_LV2_HA5/X_XOR/N002_XCSA/X_LV2_HA5/X_xor/M3_g
+ N_GND_XCSA/X_LV2_HA5/X_xor/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA5/M14 N_XCSA/LV2_C[8]_XCSA/X_LV2_HA5/M14_d
+ N_XCSA/X_LV2_HA5/N001_XCSA/X_LV2_HA5/M14_g N_GND_XCSA/X_LV2_HA5/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa17/Xyb3/M37 N_XADDER/XA17/XYB3/N008_XADDER/Xa17/Xyb3/M37_d
+ N_XADDER/XA17/T1_XADDER/Xa17/Xyb3/M37_g N_GND_XADDER/Xa17/Xyb3/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd29/M8 N_X02/XD29/N3_X02/xd29/M8_d N_CLK_X02/xd29/M8_g
+ N_X02/XD29/P003_X02/xd29/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa76/M2 N_XADDER/XA76/N002_XADDER/Xa76/M2_d
+ N_XADDER/GX5[0]_XADDER/Xa76/M2_g N_XADDER/P6_XADDER/Xa76/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA3/M26 N_XCSA/LV1_C[8]_XCSA/X_LV1_FA3/M26_d
+ N_XCSA/X_LV1_FA3/_COUT_XCSA/X_LV1_FA3/M26_g N_GND_XCSA/X_LV1_FA3/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa08/Xrb2/M3 N_XADDER/P7_XADDER/Xa08/Xrb2/M3_d
+ N_XADDER/XA08/XRB2/N002_XADDER/Xa08/Xrb2/M3_g N_GND_XADDER/Xa08/Xrb2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel23/M13 N_PP2[3]_XBOOTH/Xsel23/M13_d
+ N_XBOOTH/XSEL23/N004_XBOOTH/Xsel23/M13_g N_GND_XBOOTH/Xsel23/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel13/M13 N_PP1[3]_XBOOTH/Xsel13/M13_d
+ N_XBOOTH/XSEL13/N004_XBOOTH/Xsel13/M13_g N_GND_XBOOTH/Xsel13/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel03/M13 N_PP0[3]_XBOOTH/Xsel03/M13_d
+ N_XBOOTH/XSEL03/N004_XBOOTH/Xsel03/M13_g N_GND_XBOOTH/Xsel03/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mX02/xd29/M9 N_X02/XD29/P003_X02/xd29/M9_d N_X02/XD29/N1_X02/xd29/M9_g
+ N_GND_X02/xd29/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.76e-13 PD=2.8e-07 PS=8e-07
mXADDER/Xa17/Xyb3/M38 N_XADDER/XA17/XYB3/N008_XADDER/Xa17/Xyb3/M38_d
+ N_XADDER/G7_XADDER/Xa17/Xyb3/M38_g N_GND_XADDER/Xa17/Xyb3/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa5/M8 N_XCSA/XDFFA5/N3_XCSA/Xdffa5/M8_d N_CLK_XCSA/Xdffa5/M8_g
+ N_XCSA/XDFFA5/P003_XCSA/Xdffa5/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa18/M8 N_XCSA/XDFFA18/N3_XCSA/Xdffa18/M8_d N_CLK_XCSA/Xdffa18/M8_g
+ N_XCSA/XDFFA18/P003_XCSA/Xdffa18/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV1_FA3/M25 N_XCSA/LV1_S[7]_XCSA/X_LV1_FA3/M25_d
+ N_XCSA/X_LV1_FA3/_SUM_XCSA/X_LV1_FA3/M25_g N_GND_XCSA/X_LV1_FA3/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA4/M25 N_XCSA/LV3_S[6]_XCSA/X_LV3_FA4/M25_d
+ N_XCSA/X_LV3_FA4/_SUM_XCSA/X_LV3_FA4/M25_g N_GND_XCSA/X_LV3_FA4/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa66/Xao1/Xand1/M16 N_XADDER/XA66/OUT1_XADDER/Xa66/Xao1/Xand1/M16_d
+ N_XADDER/XA66/XAO1/N003_XADDER/Xa66/Xao1/Xand1/M16_g
+ N_GND_XADDER/Xa66/Xao1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa5/M9 N_XCSA/XDFFA5/P003_XCSA/Xdffa5/M9_d
+ N_XCSA/XDFFA5/N1_XCSA/Xdffa5/M9_g N_GND_XCSA/Xdffa5/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/Xdffa18/M9 N_XCSA/XDFFA18/P003_XCSA/Xdffa18/M9_d
+ N_XCSA/XDFFA18/N1_XCSA/Xdffa18/M9_g N_GND_XCSA/Xdffa18/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mX02/xd29/M11 N_OUT[8]_X02/xd29/M11_d N_X02/XD29/N3_X02/xd29/M11_g
+ N_GND_X02/xd29/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXADDER/Xa08/Xrb2/M1 N_XADDER/XA08/XRB2/N002_XADDER/Xa08/Xrb2/M1_d
+ N_C[7]_XADDER/Xa08/Xrb2/M1_g N_S[7]_XADDER/Xa08/Xrb2/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA4/M26 N_XCSA/LV3_C[7]_XCSA/X_LV3_FA4/M26_d
+ N_XCSA/X_LV3_FA4/_COUT_XCSA/X_LV3_FA4/M26_g N_GND_XCSA/X_LV3_FA4/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa78/M3 N_OUT1[8]_XADDER/Xa78/M3_d N_XADDER/XA78/N002_XADDER/Xa78/M3_g
+ N_GND_XADDER/Xa78/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa17/Xyb3/Xor1/M16 N_XADDER/GG7_XADDER/Xa17/Xyb3/Xor1/M16_d
+ N_XADDER/XA17/XYB3/N008_XADDER/Xa17/Xyb3/Xor1/M16_g
+ N_GND_XADDER/Xa17/Xyb3/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa5/M11 N_C[6]_XCSA/Xdffa5/M11_d N_XCSA/XDFFA5/N3_XCSA/Xdffa5/M11_g
+ N_GND_XCSA/Xdffa5/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/Xdffa18/M11 N_S[6]_XCSA/Xdffa18/M11_d N_XCSA/XDFFA18/N3_XCSA/Xdffa18/M11_g
+ N_GND_XCSA/Xdffa18/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/X_LV3_FA4/M21 N_XCSA/X_LV3_FA4/_SUM_XCSA/X_LV3_FA4/M21_d
+ N_XCSA/X_LV3_FA4/_COUT_XCSA/X_LV3_FA4/M21_g
+ N_XCSA/X_LV3_FA4/N004_XCSA/X_LV3_FA4/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXADDER/Xa08/Xrb2/M2 N_XADDER/XA08/XRB2/N002_XADDER/Xa08/Xrb2/M2_d
+ N_S[7]_XADDER/Xa08/Xrb2/M2_g N_C[7]_XADDER/Xa08/Xrb2/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXADDER/Xa66/Xao2/M37 N_XADDER/XA66/XAO2/N008_XADDER/Xa66/Xao2/M37_d
+ N_XADDER/XA66/OUT1_XADDER/Xa66/Xao2/M37_g N_GND_XADDER/Xa66/Xao2/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel24/M2 N_noxref_2225_XBOOTH/Xsel24/M2_d
+ N_XBOOTH/B_D[3]_XBOOTH/Xsel24/M2_g N_GND_XBOOTH/Xsel24/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel14/M2 N_noxref_2226_XBOOTH/Xsel14/M2_d
+ N_XBOOTH/B_D[3]_XBOOTH/Xsel14/M2_g N_GND_XBOOTH/Xsel14/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel04/M2 N_noxref_2227_XBOOTH/Xsel04/M2_d
+ N_XBOOTH/B_D[3]_XBOOTH/Xsel04/M2_g N_GND_XBOOTH/Xsel04/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mX02/xd210/M3 N_X02/XD210/N0_X02/xd210/M3_d N_OUT1[9]_X02/xd210/M3_g
+ N_GND_X02/xd210/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA4/M19 N_XCSA/X_LV1_FA4/N004_XCSA/X_LV1_FA4/M19_d
+ N_PP0[6]_XCSA/X_LV1_FA4/M19_g N_GND_XCSA/X_LV1_FA4/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA4/M24 N_XCSA/X_LV1_FA4/P006_XCSA/X_LV1_FA4/M24_d
+ N_PP0[6]_XCSA/X_LV1_FA4/M24_g N_GND_XCSA/X_LV1_FA4/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA4/M14 N_XCSA/X_LV1_FA4/P004_XCSA/X_LV1_FA4/M14_d
+ N_PP0[6]_XCSA/X_LV1_FA4/M14_g N_GND_XCSA/X_LV1_FA4/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA4/M16 N_XCSA/X_LV1_FA4/N003_XCSA/X_LV1_FA4/M16_d
+ N_PP0[6]_XCSA/X_LV1_FA4/M16_g N_GND_XCSA/X_LV1_FA4/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA4/M18 N_XCSA/X_LV3_FA4/N004_XCSA/X_LV3_FA4/M18_d
+ N_CACC[6]_XCSA/X_LV3_FA4/M18_g N_GND_XCSA/X_LV3_FA4/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA4/M22 N_XCSA/X_LV3_FA4/_SUM_XCSA/X_LV3_FA4/M22_d
+ N_CACC[6]_XCSA/X_LV3_FA4/M22_g N_XCSA/X_LV3_FA4/P005_XCSA/X_LV3_FA4/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV3_FA4/M15 N_XCSA/X_LV3_FA4/_COUT_XCSA/X_LV3_FA4/M15_d
+ N_CACC[6]_XCSA/X_LV3_FA4/M15_g N_XCSA/X_LV3_FA4/N003_XCSA/X_LV3_FA4/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXADDER/Xa66/Xao2/M38 N_XADDER/XA66/XAO2/N008_XADDER/Xa66/Xao2/M38_d
+ N_XADDER/G6_XADDER/Xa66/Xao2/M38_g N_GND_XADDER/Xa66/Xao2/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV2_HA6/X_xor/M2 N_XCSA/X_LV2_HA6/X_XOR/N002_XCSA/X_LV2_HA6/X_xor/M2_d
+ N_XCSA/LV1_C[8]_XCSA/X_LV2_HA6/X_xor/M2_g
+ N_XCSA/LV1_S[8]_XCSA/X_LV2_HA6/X_xor/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13 PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA6/M11 N_XCSA/X_LV2_HA6/P001_XCSA/X_LV2_HA6/M11_d
+ N_XCSA/LV1_C[8]_XCSA/X_LV2_HA6/M11_g N_GND_XCSA/X_LV2_HA6/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXBOOTH/Xsel24/M1 N_XBOOTH/XSEL24/N002_XBOOTH/Xsel24/M1_d
+ N_XBOOTH/D2_XBOOTH/Xsel24/M1_g N_noxref_2225_XBOOTH/Xsel24/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel14/M1 N_XBOOTH/XSEL14/N002_XBOOTH/Xsel14/M1_d
+ N_XBOOTH/D1_XBOOTH/Xsel14/M1_g N_noxref_2226_XBOOTH/Xsel14/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel04/M1 N_XBOOTH/XSEL04/N002_XBOOTH/Xsel04/M1_d
+ N_XBOOTH/D0_XBOOTH/Xsel04/M1_g N_noxref_2227_XBOOTH/Xsel04/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xdffb4/M3 N_XBOOTH/XDFFB4/N0_XBOOTH/Xdffb4/M3_d
+ N_B[4]_XBOOTH/Xdffb4/M3_g N_GND_XBOOTH/Xdffb4/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa6/M3 N_XCSA/XDFFA6/N0_XCSA/Xdffa6/M3_d
+ N_XCSA/LV3_C[7]_XCSA/Xdffa6/M3_g N_GND_XCSA/Xdffa6/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa19/M3 N_XCSA/XDFFA19/N0_XCSA/Xdffa19/M3_d
+ N_XCSA/LV3_S[7]_XCSA/Xdffa19/M3_g N_GND_XCSA/Xdffa19/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd210/M6 N_X02/XD210/P002_X02/xd210/M6_d N_CLK_X02/xd210/M6_g
+ N_GND_X02/xd210/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/X_LV1_FA4/M20 N_XCSA/X_LV1_FA4/N004_XCSA/X_LV1_FA4/M20_d
+ N_PP1[6]_XCSA/X_LV1_FA4/M20_g N_GND_XCSA/X_LV1_FA4/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV1_FA4/M23 N_XCSA/X_LV1_FA4/P005_XCSA/X_LV1_FA4/M23_d
+ N_PP1[6]_XCSA/X_LV1_FA4/M23_g N_XCSA/X_LV1_FA4/P006_XCSA/X_LV1_FA4/M23_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA4/M13 N_XCSA/X_LV1_FA4/_COUT_XCSA/X_LV1_FA4/M13_d
+ N_PP1[6]_XCSA/X_LV1_FA4/M13_g N_XCSA/X_LV1_FA4/P004_XCSA/X_LV1_FA4/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA4/M17 N_XCSA/X_LV1_FA4/N003_XCSA/X_LV1_FA4/M17_d
+ N_PP1[6]_XCSA/X_LV1_FA4/M17_g N_GND_XCSA/X_LV1_FA4/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXADDER/Xa78/M1 N_XADDER/XA78/N002_XADDER/Xa78/M1_d N_XADDER/P8_XADDER/Xa78/M1_g
+ N_XADDER/GOUT7_XADDER/Xa78/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=2.332e-13 PD=5.4e-07 PS=1.5e-06
mXCSA/X_LV3_FA4/M20 N_XCSA/X_LV3_FA4/N004_XCSA/X_LV3_FA4/M20_d
+ N_XCSA/LV2_S[6]_XCSA/X_LV3_FA4/M20_g N_GND_XCSA/X_LV3_FA4/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA4/M23 N_XCSA/X_LV3_FA4/P005_XCSA/X_LV3_FA4/M23_d
+ N_XCSA/LV2_S[6]_XCSA/X_LV3_FA4/M23_g
+ N_XCSA/X_LV3_FA4/P006_XCSA/X_LV3_FA4/M23_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA4/M13 N_XCSA/X_LV3_FA4/_COUT_XCSA/X_LV3_FA4/M13_d
+ N_XCSA/LV2_S[6]_XCSA/X_LV3_FA4/M13_g
+ N_XCSA/X_LV3_FA4/P004_XCSA/X_LV3_FA4/M13_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA4/M17 N_XCSA/X_LV3_FA4/N003_XCSA/X_LV3_FA4/M17_d
+ N_XCSA/LV2_S[6]_XCSA/X_LV3_FA4/M17_g N_GND_XCSA/X_LV3_FA4/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXADDER/Xa77/M2 N_XADDER/XA77/N002_XADDER/Xa77/M2_d
+ N_XADDER/GX6[2]_XADDER/Xa77/M2_g N_XADDER/P7_XADDER/Xa77/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa08/Xrb1/M10 N_XADDER/XA08/XRB1/N004_XADDER/Xa08/Xrb1/M10_d
+ N_S[7]_XADDER/Xa08/Xrb1/M10_g N_GND_XADDER/Xa08/Xrb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXCSA/X_LV2_HA6/X_xor/M1 N_XCSA/X_LV2_HA6/X_XOR/N002_XCSA/X_LV2_HA6/X_xor/M1_d
+ N_XCSA/LV1_S[8]_XCSA/X_LV2_HA6/X_xor/M1_g
+ N_XCSA/LV1_C[8]_XCSA/X_LV2_HA6/X_xor/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_HA6/M12 N_XCSA/X_LV2_HA6/N001_XCSA/X_LV2_HA6/M12_d
+ N_XCSA/LV1_S[8]_XCSA/X_LV2_HA6/M12_g
+ N_XCSA/X_LV2_HA6/P001_XCSA/X_LV2_HA6/M12_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mX02/xd210/M5 N_X02/XD210/N1_X02/xd210/M5_d N_X02/XD210/N0_X02/xd210/M5_g
+ N_X02/XD210/P002_X02/xd210/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel24/M3 N_XBOOTH/XSEL24/N002_XBOOTH/Xsel24/M3_d
+ N_XBOOTH/S2_XBOOTH/Xsel24/M3_g N_noxref_2237_XBOOTH/Xsel24/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel14/M3 N_XBOOTH/XSEL14/N002_XBOOTH/Xsel14/M3_d
+ N_XBOOTH/S1_XBOOTH/Xsel14/M3_g N_noxref_2238_XBOOTH/Xsel14/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel04/M3 N_XBOOTH/XSEL04/N002_XBOOTH/Xsel04/M3_d
+ N_XBOOTH/S0_XBOOTH/Xsel04/M3_g N_noxref_2239_XBOOTH/Xsel04/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xdffb4/M6 N_XBOOTH/XDFFB4/P002_XBOOTH/Xdffb4/M6_d
+ N_CLK_XBOOTH/Xdffb4/M6_g N_GND_XBOOTH/Xdffb4/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXCSA/Xdffa6/M6 N_XCSA/XDFFA6/P002_XCSA/Xdffa6/M6_d N_CLK_XCSA/Xdffa6/M6_g
+ N_GND_XCSA/Xdffa6/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/Xdffa19/M6 N_XCSA/XDFFA19/P002_XCSA/Xdffa19/M6_d N_CLK_XCSA/Xdffa19/M6_g
+ N_GND_XCSA/Xdffa19/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXADDER/Xa08/Xrb1/M9 N_XADDER/XA08/XRB1/N003_XADDER/Xa08/Xrb1/M9_d
+ N_C[7]_XADDER/Xa08/Xrb1/M9_g N_XADDER/XA08/XRB1/N004_XADDER/Xa08/Xrb1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14
+ PD=1.44e-06 PS=2.8e-07
mXCSA/X_LV1_FA4/M18 N_XCSA/X_LV1_FA4/N004_XCSA/X_LV1_FA4/M18_d
+ N_PP2[4]_XCSA/X_LV1_FA4/M18_g N_GND_XCSA/X_LV1_FA4/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV1_FA4/M22 N_XCSA/X_LV1_FA4/_SUM_XCSA/X_LV1_FA4/M22_d
+ N_PP2[4]_XCSA/X_LV1_FA4/M22_g N_XCSA/X_LV1_FA4/P005_XCSA/X_LV1_FA4/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV1_FA4/M15 N_XCSA/X_LV1_FA4/_COUT_XCSA/X_LV1_FA4/M15_d
+ N_PP2[4]_XCSA/X_LV1_FA4/M15_g N_XCSA/X_LV1_FA4/N003_XCSA/X_LV1_FA4/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXADDER/Xa66/Xao2/Xor1/M16 N_XADDER/GX6[2]_XADDER/Xa66/Xao2/Xor1/M16_d
+ N_XADDER/XA66/XAO2/N008_XADDER/Xa66/Xao2/Xor1/M16_g
+ N_GND_XADDER/Xa66/Xao2/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa78/M2 N_XADDER/XA78/N002_XADDER/Xa78/M2_d
+ N_XADDER/GOUT7_XADDER/Xa78/M2_g N_XADDER/P8_XADDER/Xa78/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xdffb4/M5 N_XBOOTH/XDFFB4/N1_XBOOTH/Xdffb4/M5_d
+ N_XBOOTH/XDFFB4/N0_XBOOTH/Xdffb4/M5_g N_XBOOTH/XDFFB4/P002_XBOOTH/Xdffb4/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV3_FA4/M19 N_XCSA/X_LV3_FA4/N004_XCSA/X_LV3_FA4/M19_d
+ N_XCSA/LV2_C[6]_XCSA/X_LV3_FA4/M19_g N_GND_XCSA/X_LV3_FA4/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA4/M24 N_XCSA/X_LV3_FA4/P006_XCSA/X_LV3_FA4/M24_d
+ N_XCSA/LV2_C[6]_XCSA/X_LV3_FA4/M24_g N_GND_XCSA/X_LV3_FA4/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA4/M14 N_XCSA/X_LV3_FA4/P004_XCSA/X_LV3_FA4/M14_d
+ N_XCSA/LV2_C[6]_XCSA/X_LV3_FA4/M14_g N_GND_XCSA/X_LV3_FA4/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA4/M16 N_XCSA/X_LV3_FA4/N003_XCSA/X_LV3_FA4/M16_d
+ N_XCSA/LV2_C[6]_XCSA/X_LV3_FA4/M16_g N_GND_XCSA/X_LV3_FA4/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa77/M1 N_XADDER/XA77/N002_XADDER/Xa77/M1_d N_XADDER/P7_XADDER/Xa77/M1_g
+ N_XADDER/GX6[2]_XADDER/Xa77/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=2.332e-13 PD=5.4e-07 PS=1.5e-06
mXCSA/Xdffa6/M5 N_XCSA/XDFFA6/N1_XCSA/Xdffa6/M5_d
+ N_XCSA/XDFFA6/N0_XCSA/Xdffa6/M5_g N_XCSA/XDFFA6/P002_XCSA/Xdffa6/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa19/M5 N_XCSA/XDFFA19/N1_XCSA/Xdffa19/M5_d
+ N_XCSA/XDFFA19/N0_XCSA/Xdffa19/M5_g N_XCSA/XDFFA19/P002_XCSA/Xdffa19/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel24/M4 N_noxref_2237_XBOOTH/Xsel24/M4_d
+ N_XBOOTH/B_D[4]_XBOOTH/Xsel24/M4_g N_GND_XBOOTH/Xsel24/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel14/M4 N_noxref_2238_XBOOTH/Xsel14/M4_d
+ N_XBOOTH/B_D[4]_XBOOTH/Xsel14/M4_g N_GND_XBOOTH/Xsel14/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel04/M4 N_noxref_2239_XBOOTH/Xsel04/M4_d
+ N_XBOOTH/B_D[4]_XBOOTH/Xsel04/M4_g N_GND_XBOOTH/Xsel04/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXCSA/X_LV1_FA4/M21 N_XCSA/X_LV1_FA4/_SUM_XCSA/X_LV1_FA4/M21_d
+ N_XCSA/X_LV1_FA4/_COUT_XCSA/X_LV1_FA4/M21_g
+ N_XCSA/X_LV1_FA4/N004_XCSA/X_LV1_FA4/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXCSA/X_LV2_HA6/X_xor/M3 N_XCSA/LV2_S[8]_XCSA/X_LV2_HA6/X_xor/M3_d
+ N_XCSA/X_LV2_HA6/X_XOR/N002_XCSA/X_LV2_HA6/X_xor/M3_g
+ N_GND_XCSA/X_LV2_HA6/X_xor/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA6/M14 N_XCSA/LV2_C[9]_XCSA/X_LV2_HA6/M14_d
+ N_XCSA/X_LV2_HA6/N001_XCSA/X_LV2_HA6/M14_g N_GND_XCSA/X_LV2_HA6/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mX02/xd210/M8 N_X02/XD210/N3_X02/xd210/M8_d N_CLK_X02/xd210/M8_g
+ N_X02/XD210/P003_X02/xd210/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel24/M5 N_XBOOTH/XSEL24/B_XBOOTH/Xsel24/M5_d
+ N_XBOOTH/XSEL24/N002_XBOOTH/Xsel24/M5_g N_GND_XBOOTH/Xsel24/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel14/M5 N_XBOOTH/XSEL14/B_XBOOTH/Xsel14/M5_d
+ N_XBOOTH/XSEL14/N002_XBOOTH/Xsel14/M5_g N_GND_XBOOTH/Xsel14/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel04/M5 N_XBOOTH/XSEL04/B_XBOOTH/Xsel04/M5_d
+ N_XBOOTH/XSEL04/N002_XBOOTH/Xsel04/M5_g N_GND_XBOOTH/Xsel04/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa08/Xrb1/Xand1/M16 N_XADDER/G7_XADDER/Xa08/Xrb1/Xand1/M16_d
+ N_XADDER/XA08/XRB1/N003_XADDER/Xa08/Xrb1/Xand1/M16_g
+ N_GND_XADDER/Xa08/Xrb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA4/M26 N_XCSA/LV1_C[9]_XCSA/X_LV1_FA4/M26_d
+ N_XCSA/X_LV1_FA4/_COUT_XCSA/X_LV1_FA4/M26_g N_GND_XCSA/X_LV1_FA4/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mX02/xd210/M9 N_X02/XD210/P003_X02/xd210/M9_d N_X02/XD210/N1_X02/xd210/M9_g
+ N_GND_X02/xd210/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.76e-13 PD=2.8e-07 PS=8e-07
mXBOOTH/Xdffb4/M8 N_XBOOTH/XDFFB4/N3_XBOOTH/Xdffb4/M8_d N_CLK_XBOOTH/Xdffb4/M8_g
+ N_XBOOTH/XDFFB4/P003_XBOOTH/Xdffb4/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV3_FA5/M25 N_XCSA/LV3_S[7]_XCSA/X_LV3_FA5/M25_d
+ N_XCSA/X_LV3_FA5/_SUM_XCSA/X_LV3_FA5/M25_g N_GND_XCSA/X_LV3_FA5/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa6/M8 N_XCSA/XDFFA6/N3_XCSA/Xdffa6/M8_d N_CLK_XCSA/Xdffa6/M8_g
+ N_XCSA/XDFFA6/P003_XCSA/Xdffa6/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa19/M8 N_XCSA/XDFFA19/N3_XCSA/Xdffa19/M8_d N_CLK_XCSA/Xdffa19/M8_g
+ N_XCSA/XDFFA19/P003_XCSA/Xdffa19/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xdffb4/M9 N_XBOOTH/XDFFB4/P003_XBOOTH/Xdffb4/M9_d
+ N_XBOOTH/XDFFB4/N1_XBOOTH/Xdffb4/M9_g N_GND_XBOOTH/Xdffb4/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXADDER/Xa77/M3 N_OUT1[7]_XADDER/Xa77/M3_d N_XADDER/XA77/N002_XADDER/Xa77/M3_g
+ N_GND_XADDER/Xa77/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa6/M9 N_XCSA/XDFFA6/P003_XCSA/Xdffa6/M9_d
+ N_XCSA/XDFFA6/N1_XCSA/Xdffa6/M9_g N_GND_XCSA/Xdffa6/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/Xdffa19/M9 N_XCSA/XDFFA19/P003_XCSA/Xdffa19/M9_d
+ N_XCSA/XDFFA19/N1_XCSA/Xdffa19/M9_g N_GND_XCSA/Xdffa19/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/X_LV1_FA4/M25 N_XCSA/LV1_S[8]_XCSA/X_LV1_FA4/M25_d
+ N_XCSA/X_LV1_FA4/_SUM_XCSA/X_LV1_FA4/M25_g N_GND_XCSA/X_LV1_FA4/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa68/Xao1/M9 N_XADDER/XA68/XAO1/N003_XADDER/Xa68/Xao1/M9_d
+ N_XADDER/GOUT7_XADDER/Xa68/Xao1/M9_g
+ N_XADDER/XA68/XAO1/N004_XADDER/Xa68/Xao1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14 PD=1.44e-06 PS=2.8e-07
mXCSA/X_LV3_FA5/M26 N_XCSA/LV3_C[8]_XCSA/X_LV3_FA5/M26_d
+ N_XCSA/X_LV3_FA5/_COUT_XCSA/X_LV3_FA5/M26_g N_GND_XCSA/X_LV3_FA5/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mX02/xd210/M11 N_OUT[9]_X02/xd210/M11_d N_X02/XD210/N3_X02/xd210/M11_g
+ N_GND_X02/xd210/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXADDER/Xa68/Xao1/M10 N_XADDER/XA68/XAO1/N004_XADDER/Xa68/Xao1/M10_d
+ N_XADDER/P8_XADDER/Xa68/Xao1/M10_g N_GND_XADDER/Xa68/Xao1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.86e-13
+ PD=2.8e-07 PS=1.74e-06
mXADDER/Xa59/Xao1/M9 N_XADDER/XA59/XAO1/N003_XADDER/Xa59/Xao1/M9_d
+ N_XADDER/GOUT7_XADDER/Xa59/Xao1/M9_g
+ N_XADDER/XA59/XAO1/N004_XADDER/Xa59/Xao1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14 PD=1.44e-06 PS=2.8e-07
mXBOOTH/Xdffb4/M11 N_XBOOTH/B_D[4]_XBOOTH/Xdffb4/M11_d
+ N_XBOOTH/XDFFB4/N3_XBOOTH/Xdffb4/M11_g N_GND_XBOOTH/Xdffb4/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXCSA/X_LV3_FA5/M21 N_XCSA/X_LV3_FA5/_SUM_XCSA/X_LV3_FA5/M21_d
+ N_XCSA/X_LV3_FA5/_COUT_XCSA/X_LV3_FA5/M21_g
+ N_XCSA/X_LV3_FA5/N004_XCSA/X_LV3_FA5/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXBOOTH/Xsel24/M12 N_XBOOTH/XSEL24/N004_XBOOTH/Xsel24/M12_d
+ N_A_D[5]_XBOOTH/Xsel24/M12_g N_XBOOTH/XSEL24/B_XBOOTH/Xsel24/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel14/M12 N_XBOOTH/XSEL14/N004_XBOOTH/Xsel14/M12_d
+ N_A_D[3]_XBOOTH/Xsel14/M12_g N_XBOOTH/XSEL14/B_XBOOTH/Xsel14/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel04/M12 N_XBOOTH/XSEL04/N004_XBOOTH/Xsel04/M12_d
+ N_A_D[1]_XBOOTH/Xsel04/M12_g N_XBOOTH/XSEL04/B_XBOOTH/Xsel04/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa09/Xrb2/M3 N_XADDER/P8_XADDER/Xa09/Xrb2/M3_d
+ N_XADDER/XA09/XRB2/N002_XADDER/Xa09/Xrb2/M3_g N_GND_XADDER/Xa09/Xrb2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa6/M11 N_C[7]_XCSA/Xdffa6/M11_d N_XCSA/XDFFA6/N3_XCSA/Xdffa6/M11_g
+ N_GND_XCSA/Xdffa6/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/Xdffa19/M11 N_S[7]_XCSA/Xdffa19/M11_d N_XCSA/XDFFA19/N3_XCSA/Xdffa19/M11_g
+ N_GND_XCSA/Xdffa19/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXADDER/Xa59/Xao1/M10 N_XADDER/XA59/XAO1/N004_XADDER/Xa59/Xao1/M10_d
+ N_XADDER/PP9_XADDER/Xa59/Xao1/M10_g N_GND_XADDER/Xa59/Xao1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.86e-13
+ PD=2.8e-07 PS=1.74e-06
mXBOOTH/Xsel24/M11 N_XBOOTH/XSEL24/N004_XBOOTH/Xsel24/M11_d
+ N_XBOOTH/XSEL24/B_XBOOTH/Xsel24/M11_g N_A_D[5]_XBOOTH/Xsel24/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel14/M11 N_XBOOTH/XSEL14/N004_XBOOTH/Xsel14/M11_d
+ N_XBOOTH/XSEL14/B_XBOOTH/Xsel14/M11_g N_A_D[3]_XBOOTH/Xsel14/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel04/M11 N_XBOOTH/XSEL04/N004_XBOOTH/Xsel04/M11_d
+ N_XBOOTH/XSEL04/B_XBOOTH/Xsel04/M11_g N_A_D[1]_XBOOTH/Xsel04/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA5/M18 N_XCSA/X_LV3_FA5/N004_XCSA/X_LV3_FA5/M18_d
+ N_CACC[7]_XCSA/X_LV3_FA5/M18_g N_GND_XCSA/X_LV3_FA5/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA5/M22 N_XCSA/X_LV3_FA5/_SUM_XCSA/X_LV3_FA5/M22_d
+ N_CACC[7]_XCSA/X_LV3_FA5/M22_g N_XCSA/X_LV3_FA5/P005_XCSA/X_LV3_FA5/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV3_FA5/M15 N_XCSA/X_LV3_FA5/_COUT_XCSA/X_LV3_FA5/M15_d
+ N_CACC[7]_XCSA/X_LV3_FA5/M15_g N_XCSA/X_LV3_FA5/N003_XCSA/X_LV3_FA5/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mX02/xd28/M3 N_X02/XD28/N0_X02/xd28/M3_d N_OUT1[7]_X02/xd28/M3_g
+ N_GND_X02/xd28/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXADDER/Xa19/Xyb1/Xand1/M16 N_XADDER/PP9_XADDER/Xa19/Xyb1/Xand1/M16_d
+ N_XADDER/XA19/XYB1/N003_XADDER/Xa19/Xyb1/Xand1/M16_g
+ N_GND_XADDER/Xa19/Xyb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa68/Xao1/Xand1/M16 N_XADDER/XA68/OUT1_XADDER/Xa68/Xao1/Xand1/M16_d
+ N_XADDER/XA68/XAO1/N003_XADDER/Xa68/Xao1/Xand1/M16_g
+ N_GND_XADDER/Xa68/Xao1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA5/M19 N_XCSA/X_LV1_FA5/N004_XCSA/X_LV1_FA5/M19_d
+ N_XCSA/PP0_INVS_XCSA/X_LV1_FA5/M19_g N_GND_XCSA/X_LV1_FA5/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA5/M24 N_XCSA/X_LV1_FA5/P006_XCSA/X_LV1_FA5/M24_d
+ N_XCSA/PP0_INVS_XCSA/X_LV1_FA5/M24_g N_GND_XCSA/X_LV1_FA5/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA5/M14 N_XCSA/X_LV1_FA5/P004_XCSA/X_LV1_FA5/M14_d
+ N_XCSA/PP0_INVS_XCSA/X_LV1_FA5/M14_g N_GND_XCSA/X_LV1_FA5/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA5/M16 N_XCSA/X_LV1_FA5/N003_XCSA/X_LV1_FA5/M16_d
+ N_XCSA/PP0_INVS_XCSA/X_LV1_FA5/M16_g N_GND_XCSA/X_LV1_FA5/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa09/Xrb2/M1 N_XADDER/XA09/XRB2/N002_XADDER/Xa09/Xrb2/M1_d
+ N_C[8]_XADDER/Xa09/Xrb2/M1_g N_S[8]_XADDER/Xa09/Xrb2/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/Xdffa7/M3 N_XCSA/XDFFA7/N0_XCSA/Xdffa7/M3_d
+ N_XCSA/LV3_C[8]_XCSA/Xdffa7/M3_g N_GND_XCSA/Xdffa7/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa20/M3 N_XCSA/XDFFA20/N0_XCSA/Xdffa20/M3_d
+ N_XCSA/LV3_S[8]_XCSA/Xdffa20/M3_g N_GND_XCSA/Xdffa20/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA5/M20 N_XCSA/X_LV3_FA5/N004_XCSA/X_LV3_FA5/M20_d
+ N_XCSA/LV2_S[7]_XCSA/X_LV3_FA5/M20_g N_GND_XCSA/X_LV3_FA5/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA5/M23 N_XCSA/X_LV3_FA5/P005_XCSA/X_LV3_FA5/M23_d
+ N_XCSA/LV2_S[7]_XCSA/X_LV3_FA5/M23_g
+ N_XCSA/X_LV3_FA5/P006_XCSA/X_LV3_FA5/M23_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA5/M13 N_XCSA/X_LV3_FA5/_COUT_XCSA/X_LV3_FA5/M13_d
+ N_XCSA/LV2_S[7]_XCSA/X_LV3_FA5/M13_g
+ N_XCSA/X_LV3_FA5/P004_XCSA/X_LV3_FA5/M13_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA5/M17 N_XCSA/X_LV3_FA5/N003_XCSA/X_LV3_FA5/M17_d
+ N_XCSA/LV2_S[7]_XCSA/X_LV3_FA5/M17_g N_GND_XCSA/X_LV3_FA5/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mX02/xd28/M6 N_X02/XD28/P002_X02/xd28/M6_d N_CLK_X02/xd28/M6_g
+ N_GND_X02/xd28/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXBOOTH/Xsel24/M13 N_PP2[4]_XBOOTH/Xsel24/M13_d
+ N_XBOOTH/XSEL24/N004_XBOOTH/Xsel24/M13_g N_GND_XBOOTH/Xsel24/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel14/M13 N_PP1[4]_XBOOTH/Xsel14/M13_d
+ N_XBOOTH/XSEL14/N004_XBOOTH/Xsel14/M13_g N_GND_XBOOTH/Xsel14/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel04/M13 N_PP0[4]_XBOOTH/Xsel04/M13_d
+ N_XBOOTH/XSEL04/N004_XBOOTH/Xsel04/M13_g N_GND_XBOOTH/Xsel04/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa59/Xao1/Xand1/M16 N_XADDER/XA59/OUT1_XADDER/Xa59/Xao1/Xand1/M16_d
+ N_XADDER/XA59/XAO1/N003_XADDER/Xa59/Xao1/Xand1/M16_g
+ N_GND_XADDER/Xa59/Xao1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA5/M20 N_XCSA/X_LV1_FA5/N004_XCSA/X_LV1_FA5/M20_d
+ N_XCSA/PP1_INVS_XCSA/X_LV1_FA5/M20_g N_GND_XCSA/X_LV1_FA5/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV1_FA5/M23 N_XCSA/X_LV1_FA5/P005_XCSA/X_LV1_FA5/M23_d
+ N_XCSA/PP1_INVS_XCSA/X_LV1_FA5/M23_g
+ N_XCSA/X_LV1_FA5/P006_XCSA/X_LV1_FA5/M23_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA5/M13 N_XCSA/X_LV1_FA5/_COUT_XCSA/X_LV1_FA5/M13_d
+ N_XCSA/PP1_INVS_XCSA/X_LV1_FA5/M13_g
+ N_XCSA/X_LV1_FA5/P004_XCSA/X_LV1_FA5/M13_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA5/M17 N_XCSA/X_LV1_FA5/N003_XCSA/X_LV1_FA5/M17_d
+ N_XCSA/PP1_INVS_XCSA/X_LV1_FA5/M17_g N_GND_XCSA/X_LV1_FA5/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV2_HA7/X_xor/M2 N_XCSA/X_LV2_HA7/X_XOR/N002_XCSA/X_LV2_HA7/X_xor/M2_d
+ N_XCSA/LV1_C[9]_XCSA/X_LV2_HA7/X_xor/M2_g
+ N_XCSA/LV1_S[9]_XCSA/X_LV2_HA7/X_xor/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13 PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA7/M11 N_XCSA/X_LV2_HA7/P001_XCSA/X_LV2_HA7/M11_d
+ N_XCSA/LV1_C[9]_XCSA/X_LV2_HA7/M11_g N_GND_XCSA/X_LV2_HA7/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mX02/xd28/M5 N_X02/XD28/N1_X02/xd28/M5_d N_X02/XD28/N0_X02/xd28/M5_g
+ N_X02/XD28/P002_X02/xd28/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa09/Xrb2/M2 N_XADDER/XA09/XRB2/N002_XADDER/Xa09/Xrb2/M2_d
+ N_S[8]_XADDER/Xa09/Xrb2/M2_g N_C[8]_XADDER/Xa09/Xrb2/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/Xdffa7/M6 N_XCSA/XDFFA7/P002_XCSA/Xdffa7/M6_d N_CLK_XCSA/Xdffa7/M6_g
+ N_GND_XCSA/Xdffa7/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/Xdffa20/M6 N_XCSA/XDFFA20/P002_XCSA/Xdffa20/M6_d N_CLK_XCSA/Xdffa20/M6_g
+ N_GND_XCSA/Xdffa20/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/X_LV3_FA5/M19 N_XCSA/X_LV3_FA5/N004_XCSA/X_LV3_FA5/M19_d
+ N_XCSA/LV2_C[7]_XCSA/X_LV3_FA5/M19_g N_GND_XCSA/X_LV3_FA5/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA5/M24 N_XCSA/X_LV3_FA5/P006_XCSA/X_LV3_FA5/M24_d
+ N_XCSA/LV2_C[7]_XCSA/X_LV3_FA5/M24_g N_GND_XCSA/X_LV3_FA5/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA5/M14 N_XCSA/X_LV3_FA5/P004_XCSA/X_LV3_FA5/M14_d
+ N_XCSA/LV2_C[7]_XCSA/X_LV3_FA5/M14_g N_GND_XCSA/X_LV3_FA5/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA5/M16 N_XCSA/X_LV3_FA5/N003_XCSA/X_LV3_FA5/M16_d
+ N_XCSA/LV2_C[7]_XCSA/X_LV3_FA5/M16_g N_GND_XCSA/X_LV3_FA5/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa19/Xyb1/M9 N_XADDER/XA19/XYB1/N003_XADDER/Xa19/Xyb1/M9_d
+ N_XADDER/P8_XADDER/Xa19/Xyb1/M9_g
+ N_XADDER/XA19/XYB1/N004_XADDER/Xa19/Xyb1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=9.24e-14 PD=1.44e-06 PS=4.2e-07
mXADDER/Xa68/Xao2/M37 N_XADDER/XA68/XAO2/N008_XADDER/Xa68/Xao2/M37_d
+ N_XADDER/XA68/OUT1_XADDER/Xa68/Xao2/M37_g N_GND_XADDER/Xa68/Xao2/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa7/M5 N_XCSA/XDFFA7/N1_XCSA/Xdffa7/M5_d
+ N_XCSA/XDFFA7/N0_XCSA/Xdffa7/M5_g N_XCSA/XDFFA7/P002_XCSA/Xdffa7/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa20/M5 N_XCSA/XDFFA20/N1_XCSA/Xdffa20/M5_d
+ N_XCSA/XDFFA20/N0_XCSA/Xdffa20/M5_g N_XCSA/XDFFA20/P002_XCSA/Xdffa20/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV2_HA7/X_xor/M1 N_XCSA/X_LV2_HA7/X_XOR/N002_XCSA/X_LV2_HA7/X_xor/M1_d
+ N_XCSA/LV1_S[9]_XCSA/X_LV2_HA7/X_xor/M1_g
+ N_XCSA/LV1_C[9]_XCSA/X_LV2_HA7/X_xor/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_HA7/M12 N_XCSA/X_LV2_HA7/N001_XCSA/X_LV2_HA7/M12_d
+ N_XCSA/LV1_S[9]_XCSA/X_LV2_HA7/M12_g
+ N_XCSA/X_LV2_HA7/P001_XCSA/X_LV2_HA7/M12_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA5/M18 N_XCSA/X_LV1_FA5/N004_XCSA/X_LV1_FA5/M18_d
+ N_PP2[5]_XCSA/X_LV1_FA5/M18_g N_GND_XCSA/X_LV1_FA5/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV1_FA5/M22 N_XCSA/X_LV1_FA5/_SUM_XCSA/X_LV1_FA5/M22_d
+ N_PP2[5]_XCSA/X_LV1_FA5/M22_g N_XCSA/X_LV1_FA5/P005_XCSA/X_LV1_FA5/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV1_FA5/M15 N_XCSA/X_LV1_FA5/_COUT_XCSA/X_LV1_FA5/M15_d
+ N_PP2[5]_XCSA/X_LV1_FA5/M15_g N_XCSA/X_LV1_FA5/N003_XCSA/X_LV1_FA5/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXADDER/Xa19/Xyb1/M10 N_XADDER/XA19/XYB1/N004_XADDER/Xa19/Xyb1/M10_d
+ N_XADDER/P9_XADDER/Xa19/Xyb1/M10_g N_GND_XADDER/Xa19/Xyb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=9.24e-14 AS=2.244e-13
+ PD=4.2e-07 PS=1.46e-06
mXADDER/Xa68/Xao2/M38 N_XADDER/XA68/XAO2/N008_XADDER/Xa68/Xao2/M38_d
+ N_XADDER/G8_XADDER/Xa68/Xao2/M38_g N_GND_XADDER/Xa68/Xao2/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa59/Xao2/M37 N_XADDER/XA59/XAO2/N008_XADDER/Xa59/Xao2/M37_d
+ N_XADDER/XA59/OUT1_XADDER/Xa59/Xao2/M37_g N_GND_XADDER/Xa59/Xao2/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd28/M8 N_X02/XD28/N3_X02/xd28/M8_d N_CLK_X02/xd28/M8_g
+ N_X02/XD28/P003_X02/xd28/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV1_FA5/M21 N_XCSA/X_LV1_FA5/_SUM_XCSA/X_LV1_FA5/M21_d
+ N_XCSA/X_LV1_FA5/_COUT_XCSA/X_LV1_FA5/M21_g
+ N_XCSA/X_LV1_FA5/N004_XCSA/X_LV1_FA5/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXCSA/X_LV3_FA6/M25 N_XCSA/LV3_S[8]_XCSA/X_LV3_FA6/M25_d
+ N_XCSA/X_LV3_FA6/_SUM_XCSA/X_LV3_FA6/M25_g N_GND_XCSA/X_LV3_FA6/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa09/Xrb1/M10 N_XADDER/XA09/XRB1/N004_XADDER/Xa09/Xrb1/M10_d
+ N_S[8]_XADDER/Xa09/Xrb1/M10_g N_GND_XADDER/Xa09/Xrb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mX02/xd28/M9 N_X02/XD28/P003_X02/xd28/M9_d N_X02/XD28/N1_X02/xd28/M9_g
+ N_GND_X02/xd28/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.76e-13 PD=2.8e-07 PS=8e-07
mXBOOTH/Xsel25/M2 N_noxref_2262_XBOOTH/Xsel25/M2_d
+ N_XBOOTH/B_D[4]_XBOOTH/Xsel25/M2_g N_GND_XBOOTH/Xsel25/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel15/M2 N_noxref_2263_XBOOTH/Xsel15/M2_d
+ N_XBOOTH/B_D[4]_XBOOTH/Xsel15/M2_g N_GND_XBOOTH/Xsel15/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel05/M2 N_noxref_2264_XBOOTH/Xsel05/M2_d
+ N_XBOOTH/B_D[4]_XBOOTH/Xsel05/M2_g N_GND_XBOOTH/Xsel05/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa59/Xao2/M38 N_XADDER/XA59/XAO2/N008_XADDER/Xa59/Xao2/M38_d
+ N_XADDER/GG9_XADDER/Xa59/Xao2/M38_g N_GND_XADDER/Xa59/Xao2/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa7/M8 N_XCSA/XDFFA7/N3_XCSA/Xdffa7/M8_d N_CLK_XCSA/Xdffa7/M8_g
+ N_XCSA/XDFFA7/P003_XCSA/Xdffa7/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa20/M8 N_XCSA/XDFFA20/N3_XCSA/Xdffa20/M8_d N_CLK_XCSA/Xdffa20/M8_g
+ N_XCSA/XDFFA20/P003_XCSA/Xdffa20/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV2_HA7/X_xor/M3 N_XCSA/LV2_S[9]_XCSA/X_LV2_HA7/X_xor/M3_d
+ N_XCSA/X_LV2_HA7/X_XOR/N002_XCSA/X_LV2_HA7/X_xor/M3_g
+ N_GND_XCSA/X_LV2_HA7/X_xor/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA7/M14 N_XCSA/LV2_C[10]_XCSA/X_LV2_HA7/M14_d
+ N_XCSA/X_LV2_HA7/N001_XCSA/X_LV2_HA7/M14_g N_GND_XCSA/X_LV2_HA7/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA5/M26 N_XCSA/LV1_C[10]_XCSA/X_LV1_FA5/M26_d
+ N_XCSA/X_LV1_FA5/_COUT_XCSA/X_LV1_FA5/M26_g N_GND_XCSA/X_LV1_FA5/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa09/Xrb1/M9 N_XADDER/XA09/XRB1/N003_XADDER/Xa09/Xrb1/M9_d
+ N_C[8]_XADDER/Xa09/Xrb1/M9_g N_XADDER/XA09/XRB1/N004_XADDER/Xa09/Xrb1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14
+ PD=1.44e-06 PS=2.8e-07
mXBOOTH/Xdffb5/M3 N_XBOOTH/XDFFB5/N0_XBOOTH/Xdffb5/M3_d
+ N_B[5]_XBOOTH/Xdffb5/M3_g N_GND_XBOOTH/Xdffb5/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA6/M26 N_XCSA/LV3_C[9]_XCSA/X_LV3_FA6/M26_d
+ N_XCSA/X_LV3_FA6/_COUT_XCSA/X_LV3_FA6/M26_g N_GND_XCSA/X_LV3_FA6/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa19/Xyb2/M10 N_XADDER/XA19/XYB2/N004_XADDER/Xa19/Xyb2/M10_d
+ N_XADDER/P9_XADDER/Xa19/Xyb2/M10_g N_GND_XADDER/Xa19/Xyb2/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXCSA/Xdffa7/M9 N_XCSA/XDFFA7/P003_XCSA/Xdffa7/M9_d
+ N_XCSA/XDFFA7/N1_XCSA/Xdffa7/M9_g N_GND_XCSA/Xdffa7/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/Xdffa20/M9 N_XCSA/XDFFA20/P003_XCSA/Xdffa20/M9_d
+ N_XCSA/XDFFA20/N1_XCSA/Xdffa20/M9_g N_GND_XCSA/Xdffa20/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXBOOTH/Xsel25/M1 N_XBOOTH/XSEL25/N002_XBOOTH/Xsel25/M1_d
+ N_XBOOTH/D2_XBOOTH/Xsel25/M1_g N_noxref_2262_XBOOTH/Xsel25/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel15/M1 N_XBOOTH/XSEL15/N002_XBOOTH/Xsel15/M1_d
+ N_XBOOTH/D1_XBOOTH/Xsel15/M1_g N_noxref_2263_XBOOTH/Xsel15/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel05/M1 N_XBOOTH/XSEL05/N002_XBOOTH/Xsel05/M1_d
+ N_XBOOTH/D0_XBOOTH/Xsel05/M1_g N_noxref_2264_XBOOTH/Xsel05/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXADDER/Xa68/Xao2/Xor1/M16 N_XADDER/GX6[3]_XADDER/Xa68/Xao2/Xor1/M16_d
+ N_XADDER/XA68/XAO2/N008_XADDER/Xa68/Xao2/Xor1/M16_g
+ N_GND_XADDER/Xa68/Xao2/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd28/M11 N_OUT[7]_X02/xd28/M11_d N_X02/XD28/N3_X02/xd28/M11_g
+ N_GND_X02/xd28/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/X_LV1_FA5/M25 N_XCSA/LV1_S[9]_XCSA/X_LV1_FA5/M25_d
+ N_XCSA/X_LV1_FA5/_SUM_XCSA/X_LV1_FA5/M25_g N_GND_XCSA/X_LV1_FA5/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xdffb5/M6 N_XBOOTH/XDFFB5/P002_XBOOTH/Xdffb5/M6_d
+ N_CLK_XBOOTH/Xdffb5/M6_g N_GND_XBOOTH/Xdffb5/M6_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.188e-13
+ PD=2.8e-07 PS=5.4e-07
mXADDER/Xa19/Xyb2/M9 N_XADDER/XA19/XYB2/N003_XADDER/Xa19/Xyb2/M9_d
+ N_XADDER/G8_XADDER/Xa19/Xyb2/M9_g
+ N_XADDER/XA19/XYB2/N004_XADDER/Xa19/Xyb2/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=6.16e-14 PD=1.74e-06 PS=2.8e-07
mXCSA/X_LV3_FA6/M21 N_XCSA/X_LV3_FA6/_SUM_XCSA/X_LV3_FA6/M21_d
+ N_XCSA/X_LV3_FA6/_COUT_XCSA/X_LV3_FA6/M21_g
+ N_XCSA/X_LV3_FA6/N004_XCSA/X_LV3_FA6/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXBOOTH/Xsel25/M3 N_XBOOTH/XSEL25/N002_XBOOTH/Xsel25/M3_d
+ N_XBOOTH/S2_XBOOTH/Xsel25/M3_g N_noxref_2269_XBOOTH/Xsel25/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel15/M3 N_XBOOTH/XSEL15/N002_XBOOTH/Xsel15/M3_d
+ N_XBOOTH/S1_XBOOTH/Xsel15/M3_g N_noxref_2270_XBOOTH/Xsel15/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel05/M3 N_XBOOTH/XSEL05/N002_XBOOTH/Xsel05/M3_d
+ N_XBOOTH/S0_XBOOTH/Xsel05/M3_g N_noxref_2271_XBOOTH/Xsel05/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xdffb5/M5 N_XBOOTH/XDFFB5/N1_XBOOTH/Xdffb5/M5_d
+ N_XBOOTH/XDFFB5/N0_XBOOTH/Xdffb5/M5_g N_XBOOTH/XDFFB5/P002_XBOOTH/Xdffb5/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa59/Xao2/Xor1/M16 N_XADDER/GX5[1]_XADDER/Xa59/Xao2/Xor1/M16_d
+ N_XADDER/XA59/XAO2/N008_XADDER/Xa59/Xao2/Xor1/M16_g
+ N_GND_XADDER/Xa59/Xao2/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa7/M11 N_C[8]_XCSA/Xdffa7/M11_d N_XCSA/XDFFA7/N3_XCSA/Xdffa7/M11_g
+ N_GND_XCSA/Xdffa7/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/Xdffa20/M11 N_S[8]_XCSA/Xdffa20/M11_d N_XCSA/XDFFA20/N3_XCSA/Xdffa20/M11_g
+ N_GND_XCSA/Xdffa20/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXADDER/Xa09/Xrb1/Xand1/M16 N_XADDER/G8_XADDER/Xa09/Xrb1/Xand1/M16_d
+ N_XADDER/XA09/XRB1/N003_XADDER/Xa09/Xrb1/Xand1/M16_g
+ N_GND_XADDER/Xa09/Xrb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA6/M18 N_XCSA/X_LV3_FA6/N004_XCSA/X_LV3_FA6/M18_d
+ N_CACC[8]_XCSA/X_LV3_FA6/M18_g N_GND_XCSA/X_LV3_FA6/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA6/M22 N_XCSA/X_LV3_FA6/_SUM_XCSA/X_LV3_FA6/M22_d
+ N_CACC[8]_XCSA/X_LV3_FA6/M22_g N_XCSA/X_LV3_FA6/P005_XCSA/X_LV3_FA6/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV3_FA6/M15 N_XCSA/X_LV3_FA6/_COUT_XCSA/X_LV3_FA6/M15_d
+ N_CACC[8]_XCSA/X_LV3_FA6/M15_g N_XCSA/X_LV3_FA6/N003_XCSA/X_LV3_FA6/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXBOOTH/Xsel25/M4 N_noxref_2269_XBOOTH/Xsel25/M4_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel25/M4_g N_GND_XBOOTH/Xsel25/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel15/M4 N_noxref_2270_XBOOTH/Xsel15/M4_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel15/M4_g N_GND_XBOOTH/Xsel15/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel05/M4 N_noxref_2271_XBOOTH/Xsel05/M4_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel05/M4_g N_GND_XBOOTH/Xsel05/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXADDER/Xa19/Xyb2/Xand1/M16 N_XADDER/XA19/T1_XADDER/Xa19/Xyb2/Xand1/M16_d
+ N_XADDER/XA19/XYB2/N003_XADDER/Xa19/Xyb2/Xand1/M16_g
+ N_GND_XADDER/Xa19/Xyb2/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa79/M2 N_XADDER/XA79/N002_XADDER/Xa79/M2_d
+ N_XADDER/GX6[3]_XADDER/Xa79/M2_g N_XADDER/P9_XADDER/Xa79/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA6/M20 N_XCSA/X_LV3_FA6/N004_XCSA/X_LV3_FA6/M20_d
+ N_XCSA/LV2_S[8]_XCSA/X_LV3_FA6/M20_g N_GND_XCSA/X_LV3_FA6/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA6/M23 N_XCSA/X_LV3_FA6/P005_XCSA/X_LV3_FA6/M23_d
+ N_XCSA/LV2_S[8]_XCSA/X_LV3_FA6/M23_g
+ N_XCSA/X_LV3_FA6/P006_XCSA/X_LV3_FA6/M23_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA6/M13 N_XCSA/X_LV3_FA6/_COUT_XCSA/X_LV3_FA6/M13_d
+ N_XCSA/LV2_S[8]_XCSA/X_LV3_FA6/M13_g
+ N_XCSA/X_LV3_FA6/P004_XCSA/X_LV3_FA6/M13_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA6/M17 N_XCSA/X_LV3_FA6/N003_XCSA/X_LV3_FA6/M17_d
+ N_XCSA/LV2_S[8]_XCSA/X_LV3_FA6/M17_g N_GND_XCSA/X_LV3_FA6/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXBOOTH/Xsel25/M5 N_XBOOTH/XSEL25/B_XBOOTH/Xsel25/M5_d
+ N_XBOOTH/XSEL25/N002_XBOOTH/Xsel25/M5_g N_GND_XBOOTH/Xsel25/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel15/M5 N_XBOOTH/XSEL15/B_XBOOTH/Xsel15/M5_d
+ N_XBOOTH/XSEL15/N002_XBOOTH/Xsel15/M5_g N_GND_XBOOTH/Xsel15/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel05/M5 N_XBOOTH/XSEL05/B_XBOOTH/Xsel05/M5_d
+ N_XBOOTH/XSEL05/N002_XBOOTH/Xsel05/M5_g N_GND_XBOOTH/Xsel05/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xdffb5/M8 N_XBOOTH/XDFFB5/N3_XBOOTH/Xdffb5/M8_d N_CLK_XBOOTH/Xdffb5/M8_g
+ N_XBOOTH/XDFFB5/P003_XBOOTH/Xdffb5/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV2_HA8/X_xor/M2 N_XCSA/X_LV2_HA8/X_XOR/N002_XCSA/X_LV2_HA8/X_xor/M2_d
+ N_XCSA/LV1_C[10]_XCSA/X_LV2_HA8/X_xor/M2_g
+ N_XCSA/LV1_S[10]_XCSA/X_LV2_HA8/X_xor/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13 PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA8/M11 N_XCSA/X_LV2_HA8/P001_XCSA/X_LV2_HA8/M11_d
+ N_XCSA/LV1_C[10]_XCSA/X_LV2_HA8/M11_g N_GND_XCSA/X_LV2_HA8/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV1_HA2/M14 N_XCSA/LV1_C[11]_XCSA/X_LV1_HA2/M14_d
+ N_XCSA/X_LV1_HA2/N001_XCSA/X_LV1_HA2/M14_g N_GND_XCSA/X_LV1_HA2/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_HA2/X_xor/M3 N_XCSA/LV1_S[10]_XCSA/X_LV1_HA2/X_xor/M3_d
+ N_XCSA/X_LV1_HA2/X_XOR/N002_XCSA/X_LV1_HA2/X_xor/M3_g
+ N_GND_XCSA/X_LV1_HA2/X_xor/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa8/M3 N_XCSA/XDFFA8/N0_XCSA/Xdffa8/M3_d
+ N_XCSA/LV3_C[9]_XCSA/Xdffa8/M3_g N_GND_XCSA/Xdffa8/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa21/M3 N_XCSA/XDFFA21/N0_XCSA/Xdffa21/M3_d
+ N_XCSA/LV3_S[9]_XCSA/Xdffa21/M3_g N_GND_XCSA/Xdffa21/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xdffb5/M9 N_XBOOTH/XDFFB5/P003_XBOOTH/Xdffb5/M9_d
+ N_XBOOTH/XDFFB5/N1_XBOOTH/Xdffb5/M9_g N_GND_XBOOTH/Xdffb5/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXADDER/Xa010/Xrb2/M3 N_XADDER/P9_XADDER/Xa010/Xrb2/M3_d
+ N_XADDER/XA010/XRB2/N002_XADDER/Xa010/Xrb2/M3_g N_GND_XADDER/Xa010/Xrb2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa79/M1 N_XADDER/XA79/N002_XADDER/Xa79/M1_d N_XADDER/P9_XADDER/Xa79/M1_g
+ N_XADDER/GX6[3]_XADDER/Xa79/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.188e-13 AS=2.332e-13 PD=5.4e-07 PS=1.5e-06
mXCSA/X_LV3_FA6/M19 N_XCSA/X_LV3_FA6/N004_XCSA/X_LV3_FA6/M19_d
+ N_XCSA/LV2_C[8]_XCSA/X_LV3_FA6/M19_g N_GND_XCSA/X_LV3_FA6/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA6/M24 N_XCSA/X_LV3_FA6/P006_XCSA/X_LV3_FA6/M24_d
+ N_XCSA/LV2_C[8]_XCSA/X_LV3_FA6/M24_g N_GND_XCSA/X_LV3_FA6/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA6/M14 N_XCSA/X_LV3_FA6/P004_XCSA/X_LV3_FA6/M14_d
+ N_XCSA/LV2_C[8]_XCSA/X_LV3_FA6/M14_g N_GND_XCSA/X_LV3_FA6/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA6/M16 N_XCSA/X_LV3_FA6/N003_XCSA/X_LV3_FA6/M16_d
+ N_XCSA/LV2_C[8]_XCSA/X_LV3_FA6/M16_g N_GND_XCSA/X_LV3_FA6/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV2_HA8/X_xor/M1 N_XCSA/X_LV2_HA8/X_XOR/N002_XCSA/X_LV2_HA8/X_xor/M1_d
+ N_XCSA/LV1_S[10]_XCSA/X_LV2_HA8/X_xor/M1_g
+ N_XCSA/LV1_C[10]_XCSA/X_LV2_HA8/X_xor/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_HA8/M12 N_XCSA/X_LV2_HA8/N001_XCSA/X_LV2_HA8/M12_d
+ N_XCSA/LV1_S[10]_XCSA/X_LV2_HA8/M12_g
+ N_XCSA/X_LV2_HA8/P001_XCSA/X_LV2_HA8/M12_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa8/M6 N_XCSA/XDFFA8/P002_XCSA/Xdffa8/M6_d N_CLK_XCSA/Xdffa8/M6_g
+ N_GND_XCSA/Xdffa8/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/Xdffa21/M6 N_XCSA/XDFFA21/P002_XCSA/Xdffa21/M6_d N_CLK_XCSA/Xdffa21/M6_g
+ N_GND_XCSA/Xdffa21/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXADDER/Xa211/Xyb1/Xand1/M16 N_XADDER/PPP11_XADDER/Xa211/Xyb1/Xand1/M16_d
+ N_XADDER/XA211/XYB1/N003_XADDER/Xa211/Xyb1/Xand1/M16_g
+ N_GND_XADDER/Xa211/Xyb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa19/Xyb3/M37 N_XADDER/XA19/XYB3/N008_XADDER/Xa19/Xyb3/M37_d
+ N_XADDER/XA19/T1_XADDER/Xa19/Xyb3/M37_g N_GND_XADDER/Xa19/Xyb3/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa8/M5 N_XCSA/XDFFA8/N1_XCSA/Xdffa8/M5_d
+ N_XCSA/XDFFA8/N0_XCSA/Xdffa8/M5_g N_XCSA/XDFFA8/P002_XCSA/Xdffa8/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa21/M5 N_XCSA/XDFFA21/N1_XCSA/Xdffa21/M5_d
+ N_XCSA/XDFFA21/N0_XCSA/Xdffa21/M5_g N_XCSA/XDFFA21/P002_XCSA/Xdffa21/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xdffb5/M11 N_XBOOTH/B_D[5]_XBOOTH/Xdffb5/M11_d
+ N_XBOOTH/XDFFB5/N3_XBOOTH/Xdffb5/M11_g N_GND_XBOOTH/Xdffb5/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXCSA/X_LV1_HA2/M12 N_XCSA/X_LV1_HA2/N001_XCSA/X_LV1_HA2/M12_d
+ N_PP2[6]_XCSA/X_LV1_HA2/M12_g N_XCSA/X_LV1_HA2/P001_XCSA/X_LV1_HA2/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_HA2/X_xor/M1 N_XCSA/X_LV1_HA2/X_XOR/N002_XCSA/X_LV1_HA2/X_xor/M1_d
+ N_PP2[6]_XCSA/X_LV1_HA2/X_xor/M1_g N_VDD_XCSA/X_LV1_HA2/X_xor/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa19/Xyb3/M38 N_XADDER/XA19/XYB3/N008_XADDER/Xa19/Xyb3/M38_d
+ N_XADDER/G9_XADDER/Xa19/Xyb3/M38_g N_GND_XADDER/Xa19/Xyb3/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel25/M12 N_XBOOTH/XSEL25/N004_XBOOTH/Xsel25/M12_d
+ N_A_D[5]_XBOOTH/Xsel25/M12_g N_XBOOTH/XSEL25/B_XBOOTH/Xsel25/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel15/M12 N_XBOOTH/XSEL15/N004_XBOOTH/Xsel15/M12_d
+ N_A_D[3]_XBOOTH/Xsel15/M12_g N_XBOOTH/XSEL15/B_XBOOTH/Xsel15/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel05/M12 N_XBOOTH/XSEL05/N004_XBOOTH/Xsel05/M12_d
+ N_A_D[1]_XBOOTH/Xsel05/M12_g N_XBOOTH/XSEL05/B_XBOOTH/Xsel05/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa010/Xrb2/M1 N_XADDER/XA010/XRB2/N002_XADDER/Xa010/Xrb2/M1_d
+ N_C[9]_XADDER/Xa010/Xrb2/M1_g N_S[9]_XADDER/Xa010/Xrb2/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA7/M25 N_XCSA/LV3_S[9]_XCSA/X_LV3_FA7/M25_d
+ N_XCSA/X_LV3_FA7/_SUM_XCSA/X_LV3_FA7/M25_g N_GND_XCSA/X_LV3_FA7/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mX02/xd211/M3 N_X02/XD211/N0_X02/xd211/M3_d N_OUT1[10]_X02/xd211/M3_g
+ N_GND_X02/xd211/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV2_HA8/X_xor/M3 N_XCSA/LV2_S[10]_XCSA/X_LV2_HA8/X_xor/M3_d
+ N_XCSA/X_LV2_HA8/X_XOR/N002_XCSA/X_LV2_HA8/X_xor/M3_g
+ N_GND_XCSA/X_LV2_HA8/X_xor/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA8/M14 N_XCSA/LV2_C[11]_XCSA/X_LV2_HA8/M14_d
+ N_XCSA/X_LV2_HA8/N001_XCSA/X_LV2_HA8/M14_g N_GND_XCSA/X_LV2_HA8/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_HA2/M11 N_XCSA/X_LV1_HA2/P001_XCSA/X_LV1_HA2/M11_d
+ N_VDD_XCSA/X_LV1_HA2/M11_g N_GND_XCSA/X_LV1_HA2/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV1_HA2/X_xor/M2 N_XCSA/X_LV1_HA2/X_XOR/N002_XCSA/X_LV1_HA2/X_xor/M2_d
+ N_VDD_XCSA/X_LV1_HA2/X_xor/M2_g N_PP2[6]_XCSA/X_LV1_HA2/X_xor/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXADDER/Xa211/Xyb1/M9 N_XADDER/XA211/XYB1/N003_XADDER/Xa211/Xyb1/M9_d
+ N_XADDER/PP9_XADDER/Xa211/Xyb1/M9_g
+ N_XADDER/XA211/XYB1/N004_XADDER/Xa211/Xyb1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b
+ N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=9.24e-14 PD=1.44e-06 PS=4.2e-07
mXADDER/Xa79/M3 N_OUT1[9]_XADDER/Xa79/M3_d N_XADDER/XA79/N002_XADDER/Xa79/M3_g
+ N_GND_XADDER/Xa79/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel25/M11 N_XBOOTH/XSEL25/N004_XBOOTH/Xsel25/M11_d
+ N_XBOOTH/XSEL25/B_XBOOTH/Xsel25/M11_g N_A_D[5]_XBOOTH/Xsel25/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel15/M11 N_XBOOTH/XSEL15/N004_XBOOTH/Xsel15/M11_d
+ N_XBOOTH/XSEL15/B_XBOOTH/Xsel15/M11_g N_A_D[3]_XBOOTH/Xsel15/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel05/M11 N_XBOOTH/XSEL05/N004_XBOOTH/Xsel05/M11_d
+ N_XBOOTH/XSEL05/B_XBOOTH/Xsel05/M11_g N_A_D[1]_XBOOTH/Xsel05/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa010/Xrb2/M2 N_XADDER/XA010/XRB2/N002_XADDER/Xa010/Xrb2/M2_d
+ N_S[9]_XADDER/Xa010/Xrb2/M2_g N_C[9]_XADDER/Xa010/Xrb2/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/Xdffa8/M8 N_XCSA/XDFFA8/N3_XCSA/Xdffa8/M8_d N_CLK_XCSA/Xdffa8/M8_g
+ N_XCSA/XDFFA8/P003_XCSA/Xdffa8/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa21/M8 N_XCSA/XDFFA21/N3_XCSA/Xdffa21/M8_d N_CLK_XCSA/Xdffa21/M8_g
+ N_XCSA/XDFFA21/P003_XCSA/Xdffa21/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mX02/xd211/M6 N_X02/XD211/P002_X02/xd211/M6_d N_CLK_X02/xd211/M6_g
+ N_GND_X02/xd211/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/X_LV3_FA7/M26 N_XCSA/LV3_C[10]_XCSA/X_LV3_FA7/M26_d
+ N_XCSA/X_LV3_FA7/_COUT_XCSA/X_LV3_FA7/M26_g N_GND_XCSA/X_LV3_FA7/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa211/Xyb1/M10 N_XADDER/XA211/XYB1/N004_XADDER/Xa211/Xyb1/M10_d
+ N_XADDER/PP11_XADDER/Xa211/Xyb1/M10_g N_GND_XADDER/Xa211/Xyb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=9.24e-14 AS=2.244e-13
+ PD=4.2e-07 PS=1.46e-06
mXCSA/Xdffa8/M9 N_XCSA/XDFFA8/P003_XCSA/Xdffa8/M9_d
+ N_XCSA/XDFFA8/N1_XCSA/Xdffa8/M9_g N_GND_XCSA/Xdffa8/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/Xdffa21/M9 N_XCSA/XDFFA21/P003_XCSA/Xdffa21/M9_d
+ N_XCSA/XDFFA21/N1_XCSA/Xdffa21/M9_g N_GND_XCSA/Xdffa21/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mX02/xd211/M5 N_X02/XD211/N1_X02/xd211/M5_d N_X02/XD211/N0_X02/xd211/M5_g
+ N_X02/XD211/P002_X02/xd211/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa19/Xyb3/Xor1/M16 N_XADDER/GG9_XADDER/Xa19/Xyb3/Xor1/M16_d
+ N_XADDER/XA19/XYB3/N008_XADDER/Xa19/Xyb3/Xor1/M16_g
+ N_GND_XADDER/Xa19/Xyb3/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA7/M21 N_XCSA/X_LV3_FA7/_SUM_XCSA/X_LV3_FA7/M21_d
+ N_XCSA/X_LV3_FA7/_COUT_XCSA/X_LV3_FA7/M21_g
+ N_XCSA/X_LV3_FA7/N004_XCSA/X_LV3_FA7/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXBOOTH/Xsel25/M13 N_PP2[5]_XBOOTH/Xsel25/M13_d
+ N_XBOOTH/XSEL25/N004_XBOOTH/Xsel25/M13_g N_GND_XBOOTH/Xsel25/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel15/M13 N_PP1[5]_XBOOTH/Xsel15/M13_d
+ N_XBOOTH/XSEL15/N004_XBOOTH/Xsel15/M13_g N_GND_XBOOTH/Xsel15/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel05/M13 N_PP0[5]_XBOOTH/Xsel05/M13_d
+ N_XBOOTH/XSEL05/N004_XBOOTH/Xsel05/M13_g N_GND_XBOOTH/Xsel05/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa8/M11 N_C[9]_XCSA/Xdffa8/M11_d N_XCSA/XDFFA8/N3_XCSA/Xdffa8/M11_g
+ N_GND_XCSA/Xdffa8/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/Xdffa21/M11 N_S[9]_XCSA/Xdffa21/M11_d N_XCSA/XDFFA21/N3_XCSA/Xdffa21/M11_g
+ N_GND_XCSA/Xdffa21/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXADDER/Xa411/Xao1/M9 N_XADDER/XA411/XAO1/N003_XADDER/Xa411/Xao1/M9_d
+ N_XADDER/GOUT7_XADDER/Xa411/Xao1/M9_g
+ N_XADDER/XA411/XAO1/N004_XADDER/Xa411/Xao1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b
+ N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14 PD=1.44e-06 PS=2.8e-07
mXCSA/X_LV3_FA7/M18 N_XCSA/X_LV3_FA7/N004_XCSA/X_LV3_FA7/M18_d
+ N_CACC[9]_XCSA/X_LV3_FA7/M18_g N_GND_XCSA/X_LV3_FA7/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA7/M22 N_XCSA/X_LV3_FA7/_SUM_XCSA/X_LV3_FA7/M22_d
+ N_CACC[9]_XCSA/X_LV3_FA7/M22_g N_XCSA/X_LV3_FA7/P005_XCSA/X_LV3_FA7/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV3_FA7/M15 N_XCSA/X_LV3_FA7/_COUT_XCSA/X_LV3_FA7/M15_d
+ N_CACC[9]_XCSA/X_LV3_FA7/M15_g N_XCSA/X_LV3_FA7/N003_XCSA/X_LV3_FA7/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXADDER/Xa010/Xrb1/M10 N_XADDER/XA010/XRB1/N004_XADDER/Xa010/Xrb1/M10_d
+ N_S[9]_XADDER/Xa010/Xrb1/M10_g N_GND_XADDER/Xa010/Xrb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXADDER/Xa211/Xyb2/M10 N_XADDER/XA211/XYB2/N004_XADDER/Xa211/Xyb2/M10_d
+ N_XADDER/PP11_XADDER/Xa211/Xyb2/M10_g N_GND_XADDER/Xa211/Xyb2/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mX02/xd211/M8 N_X02/XD211/N3_X02/xd211/M8_d N_CLK_X02/xd211/M8_g
+ N_X02/XD211/P003_X02/xd211/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa411/Xao1/M10 N_XADDER/XA411/XAO1/N004_XADDER/Xa411/Xao1/M10_d
+ N_XADDER/PPP11_XADDER/Xa411/Xao1/M10_g N_GND_XADDER/Xa411/Xao1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.86e-13
+ PD=2.8e-07 PS=1.74e-06
mXADDER/Xa010/Xrb1/M9 N_XADDER/XA010/XRB1/N003_XADDER/Xa010/Xrb1/M9_d
+ N_C[9]_XADDER/Xa010/Xrb1/M9_g N_XADDER/XA010/XRB1/N004_XADDER/Xa010/Xrb1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14
+ PD=1.44e-06 PS=2.8e-07
mXADDER/Xa211/Xyb2/M9 N_XADDER/XA211/XYB2/N003_XADDER/Xa211/Xyb2/M9_d
+ N_XADDER/GG9_XADDER/Xa211/Xyb2/M9_g
+ N_XADDER/XA211/XYB2/N004_XADDER/Xa211/Xyb2/M9_s N_GND_XADDER/Xa000/Xao1/M10_b
+ N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=6.16e-14 PD=1.74e-06 PS=2.8e-07
mXCSA/X_LV3_FA7/M20 N_XCSA/X_LV3_FA7/N004_XCSA/X_LV3_FA7/M20_d
+ N_XCSA/LV2_S[9]_XCSA/X_LV3_FA7/M20_g N_GND_XCSA/X_LV3_FA7/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA7/M23 N_XCSA/X_LV3_FA7/P005_XCSA/X_LV3_FA7/M23_d
+ N_XCSA/LV2_S[9]_XCSA/X_LV3_FA7/M23_g
+ N_XCSA/X_LV3_FA7/P006_XCSA/X_LV3_FA7/M23_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA7/M13 N_XCSA/X_LV3_FA7/_COUT_XCSA/X_LV3_FA7/M13_d
+ N_XCSA/LV2_S[9]_XCSA/X_LV3_FA7/M13_g
+ N_XCSA/X_LV3_FA7/P004_XCSA/X_LV3_FA7/M13_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA7/M17 N_XCSA/X_LV3_FA7/N003_XCSA/X_LV3_FA7/M17_d
+ N_XCSA/LV2_S[9]_XCSA/X_LV3_FA7/M17_g N_GND_XCSA/X_LV3_FA7/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXADDER/Xa610/Xao1/M9 N_XADDER/XA610/XAO1/N003_XADDER/Xa610/Xao1/M9_d
+ N_XADDER/GX5[1]_XADDER/Xa610/Xao1/M9_g
+ N_XADDER/XA610/XAO1/N004_XADDER/Xa610/Xao1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b
+ N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14 PD=1.44e-06 PS=2.8e-07
mX02/xd211/M9 N_X02/XD211/P003_X02/xd211/M9_d N_X02/XD211/N1_X02/xd211/M9_g
+ N_GND_X02/xd211/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.76e-13 PD=2.8e-07 PS=8e-07
mXCSA/X_LV2_HA0/M11 N_XCSA/X_LV2_HA0/P001_XCSA/X_LV2_HA0/M11_d
+ N_PP0[0]_XCSA/X_LV2_HA0/M11_g N_GND_XCSA/X_LV2_HA0/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA0/X_xor/M2 N_XCSA/X_LV2_HA0/X_XOR/N002_XCSA/X_LV2_HA0/X_xor/M2_d
+ N_PP0[0]_XCSA/X_LV2_HA0/X_xor/M2_g N_A_D[1]_XCSA/X_LV2_HA0/X_xor/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA9/X_xor/M2 N_XCSA/X_LV2_HA9/X_XOR/N002_XCSA/X_LV2_HA9/X_xor/M2_d
+ N_XCSA/LV1_C[11]_XCSA/X_LV2_HA9/X_xor/M2_g
+ N_XCSA/PP2_INVS_XCSA/X_LV2_HA9/X_xor/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13 PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA9/M11 N_XCSA/X_LV2_HA9/P001_XCSA/X_LV2_HA9/M11_d
+ N_XCSA/LV1_C[11]_XCSA/X_LV2_HA9/M11_g N_GND_XCSA/X_LV2_HA9/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXADDER/Xa610/Xao1/M10 N_XADDER/XA610/XAO1/N004_XADDER/Xa610/Xao1/M10_d
+ N_XADDER/P10_XADDER/Xa610/Xao1/M10_g N_GND_XADDER/Xa610/Xao1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.86e-13
+ PD=2.8e-07 PS=1.74e-06
mXCSA/Xdffa9/M3 N_XCSA/XDFFA9/N0_XCSA/Xdffa9/M3_d
+ N_XCSA/LV3_C[10]_XCSA/Xdffa9/M3_g N_GND_XCSA/Xdffa9/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa22/M3 N_XCSA/XDFFA22/N0_XCSA/Xdffa22/M3_d
+ N_XCSA/LV3_S[10]_XCSA/Xdffa22/M3_g N_GND_XCSA/Xdffa22/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA7/M19 N_XCSA/X_LV3_FA7/N004_XCSA/X_LV3_FA7/M19_d
+ N_XCSA/LV2_C[9]_XCSA/X_LV3_FA7/M19_g N_GND_XCSA/X_LV3_FA7/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA7/M24 N_XCSA/X_LV3_FA7/P006_XCSA/X_LV3_FA7/M24_d
+ N_XCSA/LV2_C[9]_XCSA/X_LV3_FA7/M24_g N_GND_XCSA/X_LV3_FA7/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA7/M14 N_XCSA/X_LV3_FA7/P004_XCSA/X_LV3_FA7/M14_d
+ N_XCSA/LV2_C[9]_XCSA/X_LV3_FA7/M14_g N_GND_XCSA/X_LV3_FA7/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA7/M16 N_XCSA/X_LV3_FA7/N003_XCSA/X_LV3_FA7/M16_d
+ N_XCSA/LV2_C[9]_XCSA/X_LV3_FA7/M16_g N_GND_XCSA/X_LV3_FA7/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel26/M2 N_XBOOTH/XSEL26/P001_XBOOTH/Xsel26/M2_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel26/M2_g N_GND_XBOOTH/Xsel26/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel16/M2 N_XBOOTH/XSEL16/P001_XBOOTH/Xsel16/M2_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel16/M2_g N_GND_XBOOTH/Xsel16/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel06/M2 N_XBOOTH/XSEL06/P001_XBOOTH/Xsel06/M2_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel06/M2_g N_GND_XBOOTH/Xsel06/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_HA0/M12 N_XCSA/X_LV2_HA0/N001_XCSA/X_LV2_HA0/M12_d
+ N_A_D[1]_XCSA/X_LV2_HA0/M12_g N_XCSA/X_LV2_HA0/P001_XCSA/X_LV2_HA0/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV2_HA0/X_xor/M1 N_XCSA/X_LV2_HA0/X_XOR/N002_XCSA/X_LV2_HA0/X_xor/M1_d
+ N_A_D[1]_XCSA/X_LV2_HA0/X_xor/M1_g N_PP0[0]_XCSA/X_LV2_HA0/X_xor/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mX02/xd211/M11 N_OUT[10]_X02/xd211/M11_d N_X02/XD211/N3_X02/xd211/M11_g
+ N_GND_X02/xd211/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/X_LV2_HA9/X_xor/M1 N_XCSA/X_LV2_HA9/X_XOR/N002_XCSA/X_LV2_HA9/X_xor/M1_d
+ N_XCSA/PP2_INVS_XCSA/X_LV2_HA9/X_xor/M1_g
+ N_XCSA/LV1_C[11]_XCSA/X_LV2_HA9/X_xor/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_HA9/M12 N_XCSA/X_LV2_HA9/N001_XCSA/X_LV2_HA9/M12_d
+ N_XCSA/PP2_INVS_XCSA/X_LV2_HA9/M12_g
+ N_XCSA/X_LV2_HA9/P001_XCSA/X_LV2_HA9/M12_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXADDER/Xa010/Xrb1/Xand1/M16 N_XADDER/G9_XADDER/Xa010/Xrb1/Xand1/M16_d
+ N_XADDER/XA010/XRB1/N003_XADDER/Xa010/Xrb1/Xand1/M16_g
+ N_GND_XADDER/Xa010/Xrb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa411/Xao1/Xand1/M16 N_XADDER/XA411/OUT1_XADDER/Xa411/Xao1/Xand1/M16_d
+ N_XADDER/XA411/XAO1/N003_XADDER/Xa411/Xao1/Xand1/M16_g
+ N_GND_XADDER/Xa411/Xao1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa9/M6 N_XCSA/XDFFA9/P002_XCSA/Xdffa9/M6_d N_CLK_XCSA/Xdffa9/M6_g
+ N_GND_XCSA/Xdffa9/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/Xdffa22/M6 N_XCSA/XDFFA22/P002_XCSA/Xdffa22/M6_d N_CLK_XCSA/Xdffa22/M6_g
+ N_GND_XCSA/Xdffa22/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXADDER/Xa211/Xyb2/Xand1/M16 N_XADDER/XA211/T1_XADDER/Xa211/Xyb2/Xand1/M16_d
+ N_XADDER/XA211/XYB2/N003_XADDER/Xa211/Xyb2/Xand1/M16_g
+ N_GND_XADDER/Xa211/Xyb2/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel26/M1 N_XBOOTH/XSEL26/N002_XBOOTH/Xsel26/M1_d
+ N_XBOOTH/D2_XBOOTH/Xsel26/M1_g N_XBOOTH/XSEL26/P001_XBOOTH/Xsel26/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel16/M1 N_XBOOTH/XSEL16/N002_XBOOTH/Xsel16/M1_d
+ N_XBOOTH/D1_XBOOTH/Xsel16/M1_g N_XBOOTH/XSEL16/P001_XBOOTH/Xsel16/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel06/M1 N_XBOOTH/XSEL06/N002_XBOOTH/Xsel06/M1_d
+ N_XBOOTH/D0_XBOOTH/Xsel06/M1_g N_XBOOTH/XSEL06/P001_XBOOTH/Xsel06/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXCSA/Xdffa9/M5 N_XCSA/XDFFA9/N1_XCSA/Xdffa9/M5_d
+ N_XCSA/XDFFA9/N0_XCSA/Xdffa9/M5_g N_XCSA/XDFFA9/P002_XCSA/Xdffa9/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa22/M5 N_XCSA/XDFFA22/N1_XCSA/Xdffa22/M5_d
+ N_XCSA/XDFFA22/N0_XCSA/Xdffa22/M5_g N_XCSA/XDFFA22/P002_XCSA/Xdffa22/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa610/Xao1/Xand1/M16 N_XADDER/XA610/OUT1_XADDER/Xa610/Xao1/Xand1/M16_d
+ N_XADDER/XA610/XAO1/N003_XADDER/Xa610/Xao1/Xand1/M16_g
+ N_GND_XADDER/Xa610/Xao1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA8/M25 N_XCSA/LV3_S[10]_XCSA/X_LV3_FA8/M25_d
+ N_XCSA/X_LV3_FA8/_SUM_XCSA/X_LV3_FA8/M25_g N_GND_XCSA/X_LV3_FA8/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel26/M3 N_XBOOTH/XSEL26/N002_XBOOTH/Xsel26/M3_d
+ N_XBOOTH/S2_XBOOTH/Xsel26/M3_g N_XBOOTH/XSEL26/P002_XBOOTH/Xsel26/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel16/M3 N_XBOOTH/XSEL16/N002_XBOOTH/Xsel16/M3_d
+ N_XBOOTH/S1_XBOOTH/Xsel16/M3_g N_XBOOTH/XSEL16/P002_XBOOTH/Xsel16/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel06/M3 N_XBOOTH/XSEL06/N002_XBOOTH/Xsel06/M3_d
+ N_XBOOTH/S0_XBOOTH/Xsel06/M3_g N_XBOOTH/XSEL06/P002_XBOOTH/Xsel06/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXCSA/X_LV2_HA0/M14 N_XCSA/LV2_C[1]_XCSA/X_LV2_HA0/M14_d
+ N_XCSA/X_LV2_HA0/N001_XCSA/X_LV2_HA0/M14_g N_GND_XCSA/X_LV2_HA0/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA0/X_xor/M3 N_XCSA/LV2_S[0]_XCSA/X_LV2_HA0/X_xor/M3_d
+ N_XCSA/X_LV2_HA0/X_XOR/N002_XCSA/X_LV2_HA0/X_xor/M3_g
+ N_GND_XCSA/X_LV2_HA0/X_xor/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA9/X_xor/M3 N_XCSA/LV2_S[11]_XCSA/X_LV2_HA9/X_xor/M3_d
+ N_XCSA/X_LV2_HA9/X_XOR/N002_XCSA/X_LV2_HA9/X_xor/M3_g
+ N_GND_XCSA/X_LV2_HA9/X_xor/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA9/M14 N_XCSA/LV2_C[12]_XCSA/X_LV2_HA9/M14_d
+ N_XCSA/X_LV2_HA9/N001_XCSA/X_LV2_HA9/M14_g N_GND_XCSA/X_LV2_HA9/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa411/Xao2/M37 N_XADDER/XA411/XAO2/N008_XADDER/Xa411/Xao2/M37_d
+ N_XADDER/XA411/OUT1_XADDER/Xa411/Xao2/M37_g N_GND_XADDER/Xa411/Xao2/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa011/Xrb2/M3 N_XADDER/P10_XADDER/Xa011/Xrb2/M3_d
+ N_XADDER/XA011/XRB2/N002_XADDER/Xa011/Xrb2/M3_g N_GND_XADDER/Xa011/Xrb2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa211/Xyb3/M37 N_XADDER/XA211/XYB3/N008_XADDER/Xa211/Xyb3/M37_d
+ N_XADDER/XA211/T1_XADDER/Xa211/Xyb3/M37_g N_GND_XADDER/Xa211/Xyb3/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel26/M4 N_XBOOTH/XSEL26/P002_XBOOTH/Xsel26/M4_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel26/M4_g N_GND_XBOOTH/Xsel26/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel16/M4 N_XBOOTH/XSEL16/P002_XBOOTH/Xsel16/M4_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel16/M4_g N_GND_XBOOTH/Xsel16/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel06/M4 N_XBOOTH/XSEL06/P002_XBOOTH/Xsel06/M4_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel06/M4_g N_GND_XBOOTH/Xsel06/M4_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXCSA/X_LV3_FA8/M26 N_XCSA/LV3_C[11]_XCSA/X_LV3_FA8/M26_d
+ N_XCSA/X_LV3_FA8/_COUT_XCSA/X_LV3_FA8/M26_g N_GND_XCSA/X_LV3_FA8/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa9/M8 N_XCSA/XDFFA9/N3_XCSA/Xdffa9/M8_d N_CLK_XCSA/Xdffa9/M8_g
+ N_XCSA/XDFFA9/P003_XCSA/Xdffa9/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa22/M8 N_XCSA/XDFFA22/N3_XCSA/Xdffa22/M8_d N_CLK_XCSA/Xdffa22/M8_g
+ N_XCSA/XDFFA22/P003_XCSA/Xdffa22/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa411/Xao2/M38 N_XADDER/XA411/XAO2/N008_XADDER/Xa411/Xao2/M38_d
+ N_XADDER/GGG11_XADDER/Xa411/Xao2/M38_g N_GND_XADDER/Xa411/Xao2/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa610/Xao2/M37 N_XADDER/XA610/XAO2/N008_XADDER/Xa610/Xao2/M37_d
+ N_XADDER/XA610/OUT1_XADDER/Xa610/Xao2/M37_g N_GND_XADDER/Xa610/Xao2/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA8/M21 N_XCSA/X_LV3_FA8/_SUM_XCSA/X_LV3_FA8/M21_d
+ N_XCSA/X_LV3_FA8/_COUT_XCSA/X_LV3_FA8/M21_g
+ N_XCSA/X_LV3_FA8/N004_XCSA/X_LV3_FA8/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXADDER/Xa211/Xyb3/M38 N_XADDER/XA211/XYB3/N008_XADDER/Xa211/Xyb3/M38_d
+ N_XADDER/GG11_XADDER/Xa211/Xyb3/M38_g N_GND_XADDER/Xa211/Xyb3/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa9/M9 N_XCSA/XDFFA9/P003_XCSA/Xdffa9/M9_d
+ N_XCSA/XDFFA9/N1_XCSA/Xdffa9/M9_g N_GND_XCSA/Xdffa9/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/Xdffa22/M9 N_XCSA/XDFFA22/P003_XCSA/Xdffa22/M9_d
+ N_XCSA/XDFFA22/N1_XCSA/Xdffa22/M9_g N_GND_XCSA/Xdffa22/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXBOOTH/Xsel26/M5 N_XBOOTH/XSEL26/B_XBOOTH/Xsel26/M5_d
+ N_XBOOTH/XSEL26/N002_XBOOTH/Xsel26/M5_g N_GND_XBOOTH/Xsel26/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel16/M5 N_XBOOTH/XSEL16/B_XBOOTH/Xsel16/M5_d
+ N_XBOOTH/XSEL16/N002_XBOOTH/Xsel16/M5_g N_GND_XBOOTH/Xsel16/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel06/M5 N_XBOOTH/XSEL06/B_XBOOTH/Xsel06/M5_d
+ N_XBOOTH/XSEL06/N002_XBOOTH/Xsel06/M5_g N_GND_XBOOTH/Xsel06/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa011/Xrb2/M1 N_XADDER/XA011/XRB2/N002_XADDER/Xa011/Xrb2/M1_d
+ N_C[10]_XADDER/Xa011/Xrb2/M1_g N_S[10]_XADDER/Xa011/Xrb2/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa610/Xao2/M38 N_XADDER/XA610/XAO2/N008_XADDER/Xa610/Xao2/M38_d
+ N_XADDER/G10_XADDER/Xa610/Xao2/M38_g N_GND_XADDER/Xa610/Xao2/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA8/M18 N_XCSA/X_LV3_FA8/N004_XCSA/X_LV3_FA8/M18_d
+ N_CACC[10]_XCSA/X_LV3_FA8/M18_g N_GND_XCSA/X_LV3_FA8/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA8/M22 N_XCSA/X_LV3_FA8/_SUM_XCSA/X_LV3_FA8/M22_d
+ N_CACC[10]_XCSA/X_LV3_FA8/M22_g N_XCSA/X_LV3_FA8/P005_XCSA/X_LV3_FA8/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV3_FA8/M15 N_XCSA/X_LV3_FA8/_COUT_XCSA/X_LV3_FA8/M15_d
+ N_CACC[10]_XCSA/X_LV3_FA8/M15_g N_XCSA/X_LV3_FA8/N003_XCSA/X_LV3_FA8/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV3_FA10/M19 N_XCSA/X_LV3_FA10/N004_XCSA/X_LV3_FA10/M19_d
+ N_XCSA/LV2_C[12]_XCSA/X_LV3_FA10/M19_g N_GND_XCSA/X_LV3_FA10/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA10/M24 N_XCSA/X_LV3_FA10/P006_XCSA/X_LV3_FA10/M24_d
+ N_XCSA/LV2_C[12]_XCSA/X_LV3_FA10/M24_g N_GND_XCSA/X_LV3_FA10/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA10/M14 N_XCSA/X_LV3_FA10/P004_XCSA/X_LV3_FA10/M14_d
+ N_XCSA/LV2_C[12]_XCSA/X_LV3_FA10/M14_g N_GND_XCSA/X_LV3_FA10/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA10/M16 N_XCSA/X_LV3_FA10/N003_XCSA/X_LV3_FA10/M16_d
+ N_XCSA/LV2_C[12]_XCSA/X_LV3_FA10/M16_g N_GND_XCSA/X_LV3_FA10/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa9/M11 N_C[10]_XCSA/Xdffa9/M11_d N_XCSA/XDFFA9/N3_XCSA/Xdffa9/M11_g
+ N_GND_XCSA/Xdffa9/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/Xdffa22/M11 N_S[10]_XCSA/Xdffa22/M11_d
+ N_XCSA/XDFFA22/N3_XCSA/Xdffa22/M11_g N_GND_XCSA/Xdffa22/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXCSA/X_LV3_FA9/M16 N_XCSA/X_LV3_FA9/N003_XCSA/X_LV3_FA9/M16_d
+ N_XCSA/LV2_C[11]_XCSA/X_LV3_FA9/M16_g N_GND_XCSA/X_LV3_FA9/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA9/M14 N_XCSA/X_LV3_FA9/P004_XCSA/X_LV3_FA9/M14_d
+ N_XCSA/LV2_C[11]_XCSA/X_LV3_FA9/M14_g N_GND_XCSA/X_LV3_FA9/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA9/M24 N_XCSA/X_LV3_FA9/P006_XCSA/X_LV3_FA9/M24_d
+ N_XCSA/LV2_C[11]_XCSA/X_LV3_FA9/M24_g N_GND_XCSA/X_LV3_FA9/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA9/M19 N_XCSA/X_LV3_FA9/N004_XCSA/X_LV3_FA9/M19_d
+ N_XCSA/LV2_C[11]_XCSA/X_LV3_FA9/M19_g N_GND_XCSA/X_LV3_FA9/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa411/Xao2/Xor1/M16 N_XADDER/FG11_XADDER/Xa411/Xao2/Xor1/M16_d
+ N_XADDER/XA411/XAO2/N008_XADDER/Xa411/Xao2/Xor1/M16_g
+ N_GND_XADDER/Xa411/Xao2/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa011/Xrb2/M2 N_XADDER/XA011/XRB2/N002_XADDER/Xa011/Xrb2/M2_d
+ N_S[10]_XADDER/Xa011/Xrb2/M2_g N_C[10]_XADDER/Xa011/Xrb2/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXADDER/Xa211/Xyb3/Xor1/M16 N_XADDER/GGG11_XADDER/Xa211/Xyb3/Xor1/M16_d
+ N_XADDER/XA211/XYB3/N008_XADDER/Xa211/Xyb3/Xor1/M16_g
+ N_GND_XADDER/Xa211/Xyb3/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA8/M20 N_XCSA/X_LV3_FA8/N004_XCSA/X_LV3_FA8/M20_d
+ N_XCSA/LV2_S[10]_XCSA/X_LV3_FA8/M20_g N_GND_XCSA/X_LV3_FA8/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA8/M23 N_XCSA/X_LV3_FA8/P005_XCSA/X_LV3_FA8/M23_d
+ N_XCSA/LV2_S[10]_XCSA/X_LV3_FA8/M23_g
+ N_XCSA/X_LV3_FA8/P006_XCSA/X_LV3_FA8/M23_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA8/M13 N_XCSA/X_LV3_FA8/_COUT_XCSA/X_LV3_FA8/M13_d
+ N_XCSA/LV2_S[10]_XCSA/X_LV3_FA8/M13_g
+ N_XCSA/X_LV3_FA8/P004_XCSA/X_LV3_FA8/M13_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA8/M17 N_XCSA/X_LV3_FA8/N003_XCSA/X_LV3_FA8/M17_d
+ N_XCSA/LV2_S[10]_XCSA/X_LV3_FA8/M17_g N_GND_XCSA/X_LV3_FA8/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA10/M20 N_XCSA/X_LV3_FA10/N004_XCSA/X_LV3_FA10/M20_d
+ N_VDD_XCSA/X_LV3_FA10/M20_g N_GND_XCSA/X_LV3_FA10/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA10/M23 N_XCSA/X_LV3_FA10/P005_XCSA/X_LV3_FA10/M23_d
+ N_VDD_XCSA/X_LV3_FA10/M23_g N_XCSA/X_LV3_FA10/P006_XCSA/X_LV3_FA10/M23_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA10/M13 N_XCSA/X_LV3_FA10/_COUT_XCSA/X_LV3_FA10/M13_d
+ N_VDD_XCSA/X_LV3_FA10/M13_g N_XCSA/X_LV3_FA10/P004_XCSA/X_LV3_FA10/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA10/M17 N_XCSA/X_LV3_FA10/N003_XCSA/X_LV3_FA10/M17_d
+ N_VDD_XCSA/X_LV3_FA10/M17_g N_GND_XCSA/X_LV3_FA10/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA9/M17 N_XCSA/X_LV3_FA9/N003_XCSA/X_LV3_FA9/M17_d
+ N_XCSA/LV2_S[11]_XCSA/X_LV3_FA9/M17_g N_GND_XCSA/X_LV3_FA9/M17_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA9/M13 N_XCSA/X_LV3_FA9/_COUT_XCSA/X_LV3_FA9/M13_d
+ N_XCSA/LV2_S[11]_XCSA/X_LV3_FA9/M13_g
+ N_XCSA/X_LV3_FA9/P004_XCSA/X_LV3_FA9/M13_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA9/M23 N_XCSA/X_LV3_FA9/P005_XCSA/X_LV3_FA9/M23_d
+ N_XCSA/LV2_S[11]_XCSA/X_LV3_FA9/M23_g
+ N_XCSA/X_LV3_FA9/P006_XCSA/X_LV3_FA9/M23_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=1.188e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA9/M20 N_XCSA/X_LV3_FA9/N004_XCSA/X_LV3_FA9/M20_d
+ N_XCSA/LV2_S[11]_XCSA/X_LV3_FA9/M20_g N_GND_XCSA/X_LV3_FA9/M20_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.298e-13
+ PD=5.4e-07 PS=5.9e-07
mXBOOTH/Xsel26/M12 N_XBOOTH/XSEL26/N004_XBOOTH/Xsel26/M12_d
+ N_A_D[5]_XBOOTH/Xsel26/M12_g N_XBOOTH/XSEL26/B_XBOOTH/Xsel26/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel16/M12 N_XBOOTH/XSEL16/N004_XBOOTH/Xsel16/M12_d
+ N_A_D[3]_XBOOTH/Xsel16/M12_g N_XBOOTH/XSEL16/B_XBOOTH/Xsel16/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel06/M12 N_XBOOTH/XSEL06/N004_XBOOTH/Xsel06/M12_d
+ N_A_D[1]_XBOOTH/Xsel06/M12_g N_XBOOTH/XSEL06/B_XBOOTH/Xsel06/M12_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa610/Xao2/Xor1/M16 N_XADDER/GX6[4]_XADDER/Xa610/Xao2/Xor1/M16_d
+ N_XADDER/XA610/XAO2/N008_XADDER/Xa610/Xao2/Xor1/M16_g
+ N_GND_XADDER/Xa610/Xao2/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd212/M3 N_X02/XD212/N0_X02/xd212/M3_d N_OUT1[11]_X02/xd212/M3_g
+ N_GND_X02/xd212/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA8/M19 N_XCSA/X_LV3_FA8/N004_XCSA/X_LV3_FA8/M19_d
+ N_XCSA/LV2_C[10]_XCSA/X_LV3_FA8/M19_g N_GND_XCSA/X_LV3_FA8/M19_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA8/M24 N_XCSA/X_LV3_FA8/P006_XCSA/X_LV3_FA8/M24_d
+ N_XCSA/LV2_C[10]_XCSA/X_LV3_FA8/M24_g N_GND_XCSA/X_LV3_FA8/M24_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA8/M14 N_XCSA/X_LV3_FA8/P004_XCSA/X_LV3_FA8/M14_d
+ N_XCSA/LV2_C[10]_XCSA/X_LV3_FA8/M14_g N_GND_XCSA/X_LV3_FA8/M14_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA8/M16 N_XCSA/X_LV3_FA8/N003_XCSA/X_LV3_FA8/M16_d
+ N_XCSA/LV2_C[10]_XCSA/X_LV3_FA8/M16_g N_GND_XCSA/X_LV3_FA8/M16_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA10/M18 N_XCSA/X_LV3_FA10/N004_XCSA/X_LV3_FA10/M18_d
+ N_CACC[11]_XCSA/X_LV3_FA10/M18_g N_GND_XCSA/X_LV3_FA10/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA10/M22 N_XCSA/X_LV3_FA10/_SUM_XCSA/X_LV3_FA10/M22_d
+ N_CACC[11]_XCSA/X_LV3_FA10/M22_g N_XCSA/X_LV3_FA10/P005_XCSA/X_LV3_FA10/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV3_FA10/M15 N_XCSA/X_LV3_FA10/_COUT_XCSA/X_LV3_FA10/M15_d
+ N_CACC[11]_XCSA/X_LV3_FA10/M15_g N_XCSA/X_LV3_FA10/N003_XCSA/X_LV3_FA10/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/Xdffa10/M3 N_XCSA/XDFFA10/N0_XCSA/Xdffa10/M3_d
+ N_XCSA/LV3_C[11]_XCSA/Xdffa10/M3_g N_GND_XCSA/Xdffa10/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa23/M3 N_XCSA/XDFFA23/N0_XCSA/Xdffa23/M3_d
+ N_XCSA/LV3_S[11]_XCSA/Xdffa23/M3_g N_GND_XCSA/Xdffa23/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA9/M15 N_XCSA/X_LV3_FA9/_COUT_XCSA/X_LV3_FA9/M15_d
+ N_CACC[11]_XCSA/X_LV3_FA9/M15_g N_XCSA/X_LV3_FA9/N003_XCSA/X_LV3_FA9/M15_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV3_FA9/M22 N_XCSA/X_LV3_FA9/_SUM_XCSA/X_LV3_FA9/M22_d
+ N_CACC[11]_XCSA/X_LV3_FA9/M22_g N_XCSA/X_LV3_FA9/P005_XCSA/X_LV3_FA9/M22_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.298e-13
+ PD=1.42e-06 PS=5.9e-07
mXCSA/X_LV3_FA9/M18 N_XCSA/X_LV3_FA9/N004_XCSA/X_LV3_FA9/M18_d
+ N_CACC[11]_XCSA/X_LV3_FA9/M18_g N_GND_XCSA/X_LV3_FA9/M18_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.408e-13 AS=1.298e-13
+ PD=6.4e-07 PS=5.9e-07
mXBOOTH/Xsel26/M11 N_XBOOTH/XSEL26/N004_XBOOTH/Xsel26/M11_d
+ N_XBOOTH/XSEL26/B_XBOOTH/Xsel26/M11_g N_A_D[5]_XBOOTH/Xsel26/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel16/M11 N_XBOOTH/XSEL16/N004_XBOOTH/Xsel16/M11_d
+ N_XBOOTH/XSEL16/B_XBOOTH/Xsel16/M11_g N_A_D[3]_XBOOTH/Xsel16/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel06/M11 N_XBOOTH/XSEL06/N004_XBOOTH/Xsel06/M11_d
+ N_XBOOTH/XSEL06/B_XBOOTH/Xsel06/M11_g N_A_D[1]_XBOOTH/Xsel06/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mX02/xd212/M6 N_X02/XD212/P002_X02/xd212/M6_d N_CLK_X02/xd212/M6_g
+ N_GND_X02/xd212/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXADDER/Xa011/Xrb1/M10 N_XADDER/XA011/XRB1/N004_XADDER/Xa011/Xrb1/M10_d
+ N_S[10]_XADDER/Xa011/Xrb1/M10_g N_GND_XADDER/Xa011/Xrb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXADDER/Xa712/M2 N_XADDER/XA712/N002_XADDER/Xa712/M2_d
+ N_XADDER/FG11_XADDER/Xa712/M2_g N_XADDER/P12_XADDER/Xa712/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/Xdffa10/M6 N_XCSA/XDFFA10/P002_XCSA/Xdffa10/M6_d N_CLK_XCSA/Xdffa10/M6_g
+ N_GND_XCSA/Xdffa10/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/Xdffa23/M6 N_XCSA/XDFFA23/P002_XCSA/Xdffa23/M6_d N_CLK_XCSA/Xdffa23/M6_g
+ N_GND_XCSA/Xdffa23/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/X_LV3_FA10/M21 N_XCSA/X_LV3_FA10/_SUM_XCSA/X_LV3_FA10/M21_d
+ N_XCSA/X_LV3_FA10/_COUT_XCSA/X_LV3_FA10/M21_g
+ N_XCSA/X_LV3_FA10/N004_XCSA/X_LV3_FA10/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mX02/xd212/M5 N_X02/XD212/N1_X02/xd212/M5_d N_X02/XD212/N0_X02/xd212/M5_g
+ N_X02/XD212/P002_X02/xd212/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa011/Xrb1/M9 N_XADDER/XA011/XRB1/N003_XADDER/Xa011/Xrb1/M9_d
+ N_C[10]_XADDER/Xa011/Xrb1/M9_g N_XADDER/XA011/XRB1/N004_XADDER/Xa011/Xrb1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14
+ PD=1.44e-06 PS=2.8e-07
mXCSA/X_LV3_FA9/M21 N_XCSA/X_LV3_FA9/_SUM_XCSA/X_LV3_FA9/M21_d
+ N_XCSA/X_LV3_FA9/_COUT_XCSA/X_LV3_FA9/M21_g
+ N_XCSA/X_LV3_FA9/N004_XCSA/X_LV3_FA9/M21_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.408e-13 PD=1.42e-06 PS=6.4e-07
mXCSA/Xdffa10/M5 N_XCSA/XDFFA10/N1_XCSA/Xdffa10/M5_d
+ N_XCSA/XDFFA10/N0_XCSA/Xdffa10/M5_g N_XCSA/XDFFA10/P002_XCSA/Xdffa10/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa23/M5 N_XCSA/XDFFA23/N1_XCSA/Xdffa23/M5_d
+ N_XCSA/XDFFA23/N0_XCSA/Xdffa23/M5_g N_XCSA/XDFFA23/P002_XCSA/Xdffa23/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel26/M13 N_PP2[6]_XBOOTH/Xsel26/M13_d
+ N_XBOOTH/XSEL26/N004_XBOOTH/Xsel26/M13_g N_GND_XBOOTH/Xsel26/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel16/M13 N_PP1[6]_XBOOTH/Xsel16/M13_d
+ N_XBOOTH/XSEL16/N004_XBOOTH/Xsel16/M13_g N_GND_XBOOTH/Xsel16/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel06/M13 N_PP0[6]_XBOOTH/Xsel06/M13_d
+ N_XBOOTH/XSEL06/N004_XBOOTH/Xsel06/M13_g N_GND_XBOOTH/Xsel06/M13_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA10/M26 N_XCSA/LV3_C[13]_XCSA/X_LV3_FA10/M26_d
+ N_XCSA/X_LV3_FA10/_COUT_XCSA/X_LV3_FA10/M26_g N_GND_XCSA/X_LV3_FA10/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa710/M3 N_OUT1[10]_XADDER/Xa710/M3_d
+ N_XADDER/XA710/N002_XADDER/Xa710/M3_g N_GND_XADDER/Xa710/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa712/M1 N_XADDER/XA712/N002_XADDER/Xa712/M1_d
+ N_XADDER/P12_XADDER/Xa712/M1_g N_XADDER/FG11_XADDER/Xa712/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.332e-13
+ PD=5.4e-07 PS=1.5e-06
mXADDER/Xa111/Xyb1/Xand1/M16 N_XADDER/PP11_XADDER/Xa111/Xyb1/Xand1/M16_d
+ N_XADDER/XA111/XYB1/N003_XADDER/Xa111/Xyb1/Xand1/M16_g
+ N_GND_XADDER/Xa111/Xyb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA9/M26 N_XCSA/LV3_C[12]_XCSA/X_LV3_FA9/M26_d
+ N_XCSA/X_LV3_FA9/_COUT_XCSA/X_LV3_FA9/M26_g N_GND_XCSA/X_LV3_FA9/M26_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA10/M25 N_XCSA/LV3_S[12]_XCSA/X_LV3_FA10/M25_d
+ N_XCSA/X_LV3_FA10/_SUM_XCSA/X_LV3_FA10/M25_g N_GND_XCSA/X_LV3_FA10/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mX02/xd212/M8 N_X02/XD212/N3_X02/xd212/M8_d N_CLK_X02/xd212/M8_g
+ N_X02/XD212/P003_X02/xd212/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa011/Xrb1/Xand1/M16 N_XADDER/G10_XADDER/Xa011/Xrb1/Xand1/M16_d
+ N_XADDER/XA011/XRB1/N003_XADDER/Xa011/Xrb1/Xand1/M16_g
+ N_GND_XADDER/Xa011/Xrb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA9/M25 N_XCSA/LV3_S[11]_XCSA/X_LV3_FA9/M25_d
+ N_XCSA/X_LV3_FA9/_SUM_XCSA/X_LV3_FA9/M25_g N_GND_XCSA/X_LV3_FA9/M25_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa10/M8 N_XCSA/XDFFA10/N3_XCSA/Xdffa10/M8_d N_CLK_XCSA/Xdffa10/M8_g
+ N_XCSA/XDFFA10/P003_XCSA/Xdffa10/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa23/M8 N_XCSA/XDFFA23/N3_XCSA/Xdffa23/M8_d N_CLK_XCSA/Xdffa23/M8_g
+ N_XCSA/XDFFA23/P003_XCSA/Xdffa23/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_inv2/mn N_XCSA/PP2_INVS_XCSA/X_inv2/mn_d N_PP2[6]_XCSA/X_inv2/mn_g
+ N_GND_XCSA/X_inv2/mn_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_inv1/mn N_XCSA/PP1_INVS_XCSA/X_inv1/mn_d N_PP1[6]_XCSA/X_inv1/mn_g
+ N_GND_XCSA/X_inv1/mn_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_inv0/mn N_XCSA/PP0_INVS_XCSA/X_inv0/mn_d N_PP0[6]_XCSA/X_inv0/mn_g
+ N_GND_XCSA/X_inv0/mn_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd212/M9 N_X02/XD212/P003_X02/xd212/M9_d N_X02/XD212/N1_X02/xd212/M9_g
+ N_GND_X02/xd212/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.76e-13 PD=2.8e-07 PS=8e-07
mXADDER/Xa111/Xyb1/M9 N_XADDER/XA111/XYB1/N003_XADDER/Xa111/Xyb1/M9_d
+ N_XADDER/P10_XADDER/Xa111/Xyb1/M9_g
+ N_XADDER/XA111/XYB1/N004_XADDER/Xa111/Xyb1/M9_s N_GND_XADDER/Xa000/Xao1/M10_b
+ N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=9.24e-14 PD=1.44e-06 PS=4.2e-07
mXCSA/Xdffa10/M9 N_XCSA/XDFFA10/P003_XCSA/Xdffa10/M9_d
+ N_XCSA/XDFFA10/N1_XCSA/Xdffa10/M9_g N_GND_XCSA/Xdffa10/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/Xdffa23/M9 N_XCSA/XDFFA23/P003_XCSA/Xdffa23/M9_d
+ N_XCSA/XDFFA23/N1_XCSA/Xdffa23/M9_g N_GND_XCSA/Xdffa23/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXADDER/Xa710/M1 N_XADDER/XA710/N002_XADDER/Xa710/M1_d
+ N_XADDER/P10_XADDER/Xa710/M1_g N_XADDER/GX5[1]_XADDER/Xa710/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.332e-13
+ PD=5.4e-07 PS=1.5e-06
mXADDER/Xa712/M3 N_OUT1[12]_XADDER/Xa712/M3_d
+ N_XADDER/XA712/N002_XADDER/Xa712/M3_g N_GND_XADDER/Xa712/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa111/Xyb1/M10 N_XADDER/XA111/XYB1/N004_XADDER/Xa111/Xyb1/M10_d
+ N_XADDER/P11_XADDER/Xa111/Xyb1/M10_g N_GND_XADDER/Xa111/Xyb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=9.24e-14 AS=2.244e-13
+ PD=4.2e-07 PS=1.46e-06
mX02/xd212/M11 N_OUT[11]_X02/xd212/M11_d N_X02/XD212/N3_X02/xd212/M11_g
+ N_GND_X02/xd212/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXADDER/Xa710/M2 N_XADDER/XA710/N002_XADDER/Xa710/M2_d
+ N_XADDER/GX5[1]_XADDER/Xa710/M2_g N_XADDER/P10_XADDER/Xa710/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/Xdffa10/M11 N_C[11]_XCSA/Xdffa10/M11_d
+ N_XCSA/XDFFA10/N3_XCSA/Xdffa10/M11_g N_GND_XCSA/Xdffa10/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXCSA/Xdffa23/M11 N_S[11]_XCSA/Xdffa23/M11_d
+ N_XCSA/XDFFA23/N3_XCSA/Xdffa23/M11_g N_GND_XCSA/Xdffa23/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXADDER/Xa012/Xrb2/M3 N_XADDER/P11_XADDER/Xa012/Xrb2/M3_d
+ N_XADDER/XA012/XRB2/N002_XADDER/Xa012/Xrb2/M3_g N_GND_XADDER/Xa012/Xrb2/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa111/Xyb2/M10 N_XADDER/XA111/XYB2/N004_XADDER/Xa111/Xyb2/M10_d
+ N_XADDER/P11_XADDER/Xa111/Xyb2/M10_g N_GND_XADDER/Xa111/Xyb2/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXADDER/Xa013/M2 N_XADDER/XA013/N002_XADDER/Xa013/M2_d N_C[12]_XADDER/Xa013/M2_g
+ N_S[12]_XADDER/Xa013/M2_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mX02/xd213/M3 N_X02/XD213/N0_X02/xd213/M3_d N_OUT1[12]_X02/xd213/M3_g
+ N_GND_X02/xd213/M3_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXADDER/Xa111/Xyb2/M9 N_XADDER/XA111/XYB2/N003_XADDER/Xa111/Xyb2/M9_d
+ N_XADDER/G10_XADDER/Xa111/Xyb2/M9_g
+ N_XADDER/XA111/XYB2/N004_XADDER/Xa111/Xyb2/M9_s N_GND_XADDER/Xa000/Xao1/M10_b
+ N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=6.16e-14 PD=1.74e-06 PS=2.8e-07
mXCSA/Xdffa11/M3 N_XCSA/XDFFA11/N0_XCSA/Xdffa11/M3_d
+ N_XCSA/LV3_C[12]_XCSA/Xdffa11/M3_g N_GND_XCSA/Xdffa11/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa24/M3 N_XCSA/XDFFA24/N0_XCSA/Xdffa24/M3_d
+ N_XCSA/LV3_S[12]_XCSA/Xdffa24/M3_g N_GND_XCSA/Xdffa24/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa012/Xrb2/M1 N_XADDER/XA012/XRB2/N002_XADDER/Xa012/Xrb2/M1_d
+ N_C[11]_XADDER/Xa012/Xrb2/M1_g N_S[11]_XADDER/Xa012/Xrb2/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa013/M1 N_XADDER/XA013/N002_XADDER/Xa013/M1_d N_S[12]_XADDER/Xa013/M1_g
+ N_C[12]_XADDER/Xa013/M1_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.332e-13 PD=5.4e-07 PS=1.5e-06
mX02/xd213/M6 N_X02/XD213/P002_X02/xd213/M6_d N_CLK_X02/xd213/M6_g
+ N_GND_X02/xd213/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXADDER/Xa711/M3 N_OUT1[11]_XADDER/Xa711/M3_d
+ N_XADDER/XA711/N002_XADDER/Xa711/M3_g N_GND_XADDER/Xa711/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa11/M6 N_XCSA/XDFFA11/P002_XCSA/Xdffa11/M6_d N_CLK_XCSA/Xdffa11/M6_g
+ N_GND_XCSA/Xdffa11/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXCSA/Xdffa24/M6 N_XCSA/XDFFA24/P002_XCSA/Xdffa24/M6_d N_CLK_XCSA/Xdffa24/M6_g
+ N_GND_XCSA/Xdffa24/M6_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.188e-13 PD=2.8e-07 PS=5.4e-07
mXADDER/Xa012/Xrb2/M2 N_XADDER/XA012/XRB2/N002_XADDER/Xa012/Xrb2/M2_d
+ N_S[11]_XADDER/Xa012/Xrb2/M2_g N_C[11]_XADDER/Xa012/Xrb2/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mX02/xd213/M5 N_X02/XD213/N1_X02/xd213/M5_d N_X02/XD213/N0_X02/xd213/M5_g
+ N_X02/XD213/P002_X02/xd213/M5_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa11/M5 N_XCSA/XDFFA11/N1_XCSA/Xdffa11/M5_d
+ N_XCSA/XDFFA11/N0_XCSA/Xdffa11/M5_g N_XCSA/XDFFA11/P002_XCSA/Xdffa11/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa24/M5 N_XCSA/XDFFA24/N1_XCSA/Xdffa24/M5_d
+ N_XCSA/XDFFA24/N0_XCSA/Xdffa24/M5_g N_XCSA/XDFFA24/P002_XCSA/Xdffa24/M5_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa111/Xyb2/Xand1/M16 N_XADDER/XA111/T1_XADDER/Xa111/Xyb2/Xand1/M16_d
+ N_XADDER/XA111/XYB2/N003_XADDER/Xa111/Xyb2/Xand1/M16_g
+ N_GND_XADDER/Xa111/Xyb2/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd213/M8 N_X02/XD213/N3_X02/xd213/M8_d N_CLK_X02/xd213/M8_g
+ N_X02/XD213/P003_X02/xd213/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa013/M3 N_XADDER/P12_XADDER/Xa013/M3_d
+ N_XADDER/XA013/N002_XADDER/Xa013/M3_g N_GND_XADDER/Xa013/M3_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa012/Xrb1/M10 N_XADDER/XA012/XRB1/N004_XADDER/Xa012/Xrb1/M10_d
+ N_S[11]_XADDER/Xa012/Xrb1/M10_g N_GND_XADDER/Xa012/Xrb1/M10_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.2e-13
+ PD=2.8e-07 PS=1.44e-06
mXADDER/Xa711/M1 N_XADDER/XA711/N002_XADDER/Xa711/M1_d
+ N_XADDER/P11_XADDER/Xa711/M1_g N_XADDER/GX6[4]_XADDER/Xa711/M1_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.332e-13
+ PD=5.4e-07 PS=1.5e-06
mXCSA/Xdffa11/M8 N_XCSA/XDFFA11/N3_XCSA/Xdffa11/M8_d N_CLK_XCSA/Xdffa11/M8_g
+ N_XCSA/XDFFA11/P003_XCSA/Xdffa11/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa24/M8 N_XCSA/XDFFA24/N3_XCSA/Xdffa24/M8_d N_CLK_XCSA/Xdffa24/M8_g
+ N_XCSA/XDFFA24/P003_XCSA/Xdffa24/M8_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mX02/xd213/M9 N_X02/XD213/P003_X02/xd213/M9_d N_X02/XD213/N1_X02/xd213/M9_g
+ N_GND_X02/xd213/M9_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=1.76e-13 PD=2.8e-07 PS=8e-07
mXADDER/Xa012/Xrb1/M9 N_XADDER/XA012/XRB1/N003_XADDER/Xa012/Xrb1/M9_d
+ N_C[11]_XADDER/Xa012/Xrb1/M9_g N_XADDER/XA012/XRB1/N004_XADDER/Xa012/Xrb1/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.2e-13 AS=6.16e-14
+ PD=1.44e-06 PS=2.8e-07
mXADDER/Xa111/Xyb3/M37 N_XADDER/XA111/XYB3/N008_XADDER/Xa111/Xyb3/M37_d
+ N_XADDER/XA111/T1_XADDER/Xa111/Xyb3/M37_g N_GND_XADDER/Xa111/Xyb3/M37_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa11/M9 N_XCSA/XDFFA11/P003_XCSA/Xdffa11/M9_d
+ N_XCSA/XDFFA11/N1_XCSA/Xdffa11/M9_g N_GND_XCSA/Xdffa11/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXCSA/Xdffa24/M9 N_XCSA/XDFFA24/P003_XCSA/Xdffa24/M9_d
+ N_XCSA/XDFFA24/N1_XCSA/Xdffa24/M9_g N_GND_XCSA/Xdffa24/M9_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=1.76e-13
+ PD=2.8e-07 PS=8e-07
mXADDER/Xa711/M2 N_XADDER/XA711/N002_XADDER/Xa711/M2_d
+ N_XADDER/GX6[4]_XADDER/Xa711/M2_g N_XADDER/P11_XADDER/Xa711/M2_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa111/Xyb3/M38 N_XADDER/XA111/XYB3/N008_XADDER/Xa111/Xyb3/M38_d
+ N_XADDER/G11_XADDER/Xa111/Xyb3/M38_g N_GND_XADDER/Xa111/Xyb3/M38_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd213/M11 N_OUT[12]_X02/xd213/M11_d N_X02/XD213/N3_X02/xd213/M11_g
+ N_GND_X02/xd213/M11_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.76e-13 PD=1.42e-06 PS=8e-07
mXCSA/Xdffa11/M11 N_C[12]_XCSA/Xdffa11/M11_d
+ N_XCSA/XDFFA11/N3_XCSA/Xdffa11/M11_g N_GND_XCSA/Xdffa11/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXCSA/Xdffa24/M11 N_S[12]_XCSA/Xdffa24/M11_d
+ N_XCSA/XDFFA24/N3_XCSA/Xdffa24/M11_g N_GND_XCSA/Xdffa24/M11_s
+ N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.76e-13
+ PD=1.42e-06 PS=8e-07
mXADDER/Xa012/Xrb1/Xand1/M16 N_XADDER/G11_XADDER/Xa012/Xrb1/Xand1/M16_d
+ N_XADDER/XA012/XRB1/N003_XADDER/Xa012/Xrb1/Xand1/M16_g
+ N_GND_XADDER/Xa012/Xrb1/Xand1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa111/Xyb3/Xor1/M16 N_XADDER/GG11_XADDER/Xa111/Xyb3/Xor1/M16_d
+ N_XADDER/XA111/XYB3/N008_XADDER/Xa111/Xyb3/Xor1/M16_g
+ N_GND_XADDER/Xa111/Xyb3/Xor1/M16_s N_GND_XADDER/Xa000/Xao1/M10_b N_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa000/Xao1/M12 N_XADDER/XA000/XAO1/N003_XADDER/Xa000/Xao1/M12_d
+ N_CIN_XADDER/Xa000/Xao1/M12_g N_VDD_XADDER/Xa000/Xao1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa01/Xrb2/M4 N_XADDER/P0_XADDER/Xa01/Xrb2/M4_d
+ N_XADDER/XA01/XRB2/N002_XADDER/Xa01/Xrb2/M4_g N_VDD_XADDER/Xa01/Xrb2/M4_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa72/M4 N_OUT1[2]_XADDER/Xa72/M4_d N_XADDER/XA72/N002_XADDER/Xa72/M4_g
+ N_VDD_XADDER/Xa72/M4_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa000/Xao1/M11 N_XADDER/XA000/XAO1/N003_XADDER/Xa000/Xao1/M11_d
+ N_XADDER/P0_XADDER/Xa000/Xao1/M11_g N_VDD_XADDER/Xa000/Xao1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mXADDER/Xa70/M6 N_XADDER/XA70/N001_XADDER/Xa70/M6_d N_XADDER/P0_XADDER/Xa70/M6_g
+ N_VDD_XADDER/Xa70/M6_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xdffa4/M1 N_XBOOTH/XDFFA4/P001_XBOOTH/Xdffa4/M1_d
+ N_A[4]_XBOOTH/Xdffa4/M1_g N_VDD_XBOOTH/Xdffa4/M1_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=7.7e-14 AS=2.695e-13 PD=2.8e-07 PS=1.53e-06
mXBOOTH/Xdffa5/M1 N_XBOOTH/XDFFA5/P001_XBOOTH/Xdffa5/M1_d
+ N_A[5]_XBOOTH/Xdffa5/M1_g N_VDD_XBOOTH/Xdffa5/M1_s N_VDD_XBOOTH/Xdffa5/M1_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=7.7e-14 AS=2.695e-13 PD=2.8e-07 PS=1.53e-06
mXBOOTH/Xdffa3/M1 N_XBOOTH/XDFFA3/P001_XBOOTH/Xdffa3/M1_d
+ N_A[3]_XBOOTH/Xdffa3/M1_g N_VDD_XBOOTH/Xdffa3/M1_s N_VDD_XBOOTH/Xdffa5/M1_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=7.7e-14 AS=2.695e-13 PD=2.8e-07 PS=1.53e-06
mXBOOTH/Xdffa2/M1 N_XBOOTH/XDFFA2/P001_XBOOTH/Xdffa2/M1_d
+ N_A[2]_XBOOTH/Xdffa2/M1_g N_VDD_XBOOTH/Xdffa2/M1_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=7.7e-14 AS=2.695e-13 PD=2.8e-07 PS=1.53e-06
mXBOOTH/Xdffa0/M1 N_XBOOTH/XDFFA0/P001_XBOOTH/Xdffa0/M1_d
+ N_A[0]_XBOOTH/Xdffa0/M1_g N_VDD_XBOOTH/Xdffa0/M1_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=7.7e-14 AS=2.695e-13 PD=2.8e-07 PS=1.53e-06
mXBOOTH/Xdffa1/M1 N_XBOOTH/XDFFA1/P001_XBOOTH/Xdffa1/M1_d
+ N_A[1]_XBOOTH/Xdffa1/M1_g N_VDD_XBOOTH/Xdffa1/M1_s N_VDD_XBOOTH/Xdffa1/M1_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=7.7e-14 AS=2.695e-13 PD=2.8e-07 PS=1.53e-06
mXADDER/Xa70/M5 N_XADDER/XA70/N002_XADDER/Xa70/M5_d N_CIN_XADDER/Xa70/M5_g
+ N_XADDER/XA70/N001_XADDER/Xa70/M5_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=4.444e-13 AS=6.16e-14 PD=2.46e-06 PS=2.8e-07
mXBOOTH/Xdffa4/M2 N_XBOOTH/XDFFA4/N0_XBOOTH/Xdffa4/M2_d N_CLK_XBOOTH/Xdffa4/M2_g
+ N_XBOOTH/XDFFA4/P001_XBOOTH/Xdffa4/M2_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=7.7e-14 PD=1.53e-06 PS=2.8e-07
mXBOOTH/Xdffa5/M2 N_XBOOTH/XDFFA5/N0_XBOOTH/Xdffa5/M2_d N_CLK_XBOOTH/Xdffa5/M2_g
+ N_XBOOTH/XDFFA5/P001_XBOOTH/Xdffa5/M2_s N_VDD_XBOOTH/Xdffa5/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=7.7e-14 PD=1.53e-06 PS=2.8e-07
mXBOOTH/Xdffa3/M2 N_XBOOTH/XDFFA3/N0_XBOOTH/Xdffa3/M2_d N_CLK_XBOOTH/Xdffa3/M2_g
+ N_XBOOTH/XDFFA3/P001_XBOOTH/Xdffa3/M2_s N_VDD_XBOOTH/Xdffa5/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=7.7e-14 PD=1.53e-06 PS=2.8e-07
mXBOOTH/Xdffa2/M2 N_XBOOTH/XDFFA2/N0_XBOOTH/Xdffa2/M2_d N_CLK_XBOOTH/Xdffa2/M2_g
+ N_XBOOTH/XDFFA2/P001_XBOOTH/Xdffa2/M2_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=7.7e-14 PD=1.53e-06 PS=2.8e-07
mXBOOTH/Xdffa0/M2 N_XBOOTH/XDFFA0/N0_XBOOTH/Xdffa0/M2_d N_CLK_XBOOTH/Xdffa0/M2_g
+ N_XBOOTH/XDFFA0/P001_XBOOTH/Xdffa0/M2_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=7.7e-14 PD=1.53e-06 PS=2.8e-07
mXBOOTH/Xdffa1/M2 N_XBOOTH/XDFFA1/N0_XBOOTH/Xdffa1/M2_d N_CLK_XBOOTH/Xdffa1/M2_g
+ N_XBOOTH/XDFFA1/P001_XBOOTH/Xdffa1/M2_s N_VDD_XBOOTH/Xdffa1/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=7.7e-14 PD=1.53e-06 PS=2.8e-07
mXADDER/Xa01/Xrb2/M5 N_XADDER/XA01/XRB2/N001_XADDER/Xa01/Xrb2/M5_d
+ N_GND_XADDER/Xa01/Xrb2/M5_g N_VDD_XADDER/Xa01/Xrb2/M5_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.904e-13
+ PD=2.8e-07 PS=1.76e-06
mXADDER/Xa01/Xrb2/M6 N_XADDER/XA01/XRB2/N002_XADDER/Xa01/Xrb2/M6_d
+ N_S[0]_XADDER/Xa01/Xrb2/M6_g N_XADDER/XA01/XRB2/N001_XADDER/Xa01/Xrb2/M6_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa000/Xao1/Xand1/M15 N_VDD_XADDER/Xa000/Xao1/Xand1/M15_d
+ N_XADDER/XA000/XAO1/N003_XADDER/Xa000/Xao1/Xand1/M15_g
+ N_XADDER/XA000/OUT1_XADDER/Xa000/Xao1/Xand1/M15_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa72/M5 N_XADDER/XA72/N002_XADDER/Xa72/M5_d N_XADDER/P2_XADDER/Xa72/M5_g
+ N_XADDER/XA72/N001_XADDER/Xa72/M5_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=4.444e-13 AS=6.16e-14 PD=2.46e-06 PS=2.8e-07
mXACCXOR/X_xor1/M4 N_CACC[1]_XACCXOR/X_xor1/M4_d
+ N_XACCXOR/X_XOR1/N002_XACCXOR/X_xor1/M4_g N_VDD_XACCXOR/X_xor1/M4_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor2/M4 N_CACC[2]_XACCXOR/X_xor2/M4_d
+ N_XACCXOR/X_XOR2/N002_XACCXOR/X_xor2/M4_g N_VDD_XACCXOR/X_xor2/M4_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor4/M4 N_CACC[4]_XACCXOR/X_xor4/M4_d
+ N_XACCXOR/X_XOR4/N002_XACCXOR/X_xor4/M4_g N_VDD_XACCXOR/X_xor4/M4_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor6/M4 N_CACC[6]_XACCXOR/X_xor6/M4_d
+ N_XACCXOR/X_XOR6/N002_XACCXOR/X_xor6/M4_g N_VDD_XACCXOR/X_xor6/M4_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor8/M4 N_CACC[8]_XACCXOR/X_xor8/M4_d
+ N_XACCXOR/X_XOR8/N002_XACCXOR/X_xor8/M4_g N_VDD_XACCXOR/X_xor8/M4_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor10/M4 N_CACC[10]_XACCXOR/X_xor10/M4_d
+ N_XACCXOR/X_XOR10/N002_XACCXOR/X_xor10/M4_g N_VDD_XACCXOR/X_xor10/M4_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa72/M6 N_XADDER/XA72/N001_XADDER/Xa72/M6_d
+ N_XADDER/GG1_XADDER/Xa72/M6_g N_VDD_XADDER/Xa72/M6_s N_VDD_XADDER/Xa72/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xdffa4/M4 N_XBOOTH/XDFFA4/N1_XBOOTH/Xdffa4/M4_d N_CLK_XBOOTH/Xdffa4/M4_g
+ N_VDD_XBOOTH/Xdffa4/M4_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07
+ AD=2.695e-13 AS=1.485e-13 PD=1.53e-06 PS=5.4e-07
mXBOOTH/Xdffa5/M4 N_XBOOTH/XDFFA5/N1_XBOOTH/Xdffa5/M4_d N_CLK_XBOOTH/Xdffa5/M4_g
+ N_VDD_XBOOTH/Xdffa5/M4_s N_VDD_XBOOTH/Xdffa5/M1_b P_18_G2 L=1.8e-07 W=5.5e-07
+ AD=2.695e-13 AS=1.485e-13 PD=1.53e-06 PS=5.4e-07
mXBOOTH/Xdffa3/M4 N_XBOOTH/XDFFA3/N1_XBOOTH/Xdffa3/M4_d N_CLK_XBOOTH/Xdffa3/M4_g
+ N_VDD_XBOOTH/Xdffa3/M4_s N_VDD_XBOOTH/Xdffa5/M1_b P_18_G2 L=1.8e-07 W=5.5e-07
+ AD=2.695e-13 AS=1.485e-13 PD=1.53e-06 PS=5.4e-07
mXBOOTH/Xdffa2/M4 N_XBOOTH/XDFFA2/N1_XBOOTH/Xdffa2/M4_d N_CLK_XBOOTH/Xdffa2/M4_g
+ N_VDD_XBOOTH/Xdffa2/M4_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=5.5e-07
+ AD=2.695e-13 AS=1.485e-13 PD=1.53e-06 PS=5.4e-07
mXBOOTH/Xdffa0/M4 N_XBOOTH/XDFFA0/N1_XBOOTH/Xdffa0/M4_d N_CLK_XBOOTH/Xdffa0/M4_g
+ N_VDD_XBOOTH/Xdffa0/M4_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=5.5e-07
+ AD=2.695e-13 AS=1.485e-13 PD=1.53e-06 PS=5.4e-07
mXBOOTH/Xdffa1/M4 N_XBOOTH/XDFFA1/N1_XBOOTH/Xdffa1/M4_d N_CLK_XBOOTH/Xdffa1/M4_g
+ N_VDD_XBOOTH/Xdffa1/M4_s N_VDD_XBOOTH/Xdffa1/M1_b P_18_G2 L=1.8e-07 W=5.5e-07
+ AD=2.695e-13 AS=1.485e-13 PD=1.53e-06 PS=5.4e-07
mXADDER/Xa70/M4 N_OUT1[0]_XADDER/Xa70/M4_d N_XADDER/XA70/N002_XADDER/Xa70/M4_g
+ N_VDD_XADDER/Xa70/M4_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xdffa4/M7 N_XBOOTH/XDFFA4/N3_XBOOTH/Xdffa4/M7_d
+ N_XBOOTH/XDFFA4/N1_XBOOTH/Xdffa4/M7_g N_VDD_XBOOTH/Xdffa4/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXBOOTH/Xdffa5/M7 N_XBOOTH/XDFFA5/N3_XBOOTH/Xdffa5/M7_d
+ N_XBOOTH/XDFFA5/N1_XBOOTH/Xdffa5/M7_g N_VDD_XBOOTH/Xdffa5/M7_s
+ N_VDD_XBOOTH/Xdffa5/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXBOOTH/Xdffa3/M7 N_XBOOTH/XDFFA3/N3_XBOOTH/Xdffa3/M7_d
+ N_XBOOTH/XDFFA3/N1_XBOOTH/Xdffa3/M7_g N_VDD_XBOOTH/Xdffa3/M7_s
+ N_VDD_XBOOTH/Xdffa5/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXBOOTH/Xdffa2/M7 N_XBOOTH/XDFFA2/N3_XBOOTH/Xdffa2/M7_d
+ N_XBOOTH/XDFFA2/N1_XBOOTH/Xdffa2/M7_g N_VDD_XBOOTH/Xdffa2/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXBOOTH/Xdffa0/M7 N_XBOOTH/XDFFA0/N3_XBOOTH/Xdffa0/M7_d
+ N_XBOOTH/XDFFA0/N1_XBOOTH/Xdffa0/M7_g N_VDD_XBOOTH/Xdffa0/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXBOOTH/Xdffa1/M7 N_XBOOTH/XDFFA1/N3_XBOOTH/Xdffa1/M7_d
+ N_XBOOTH/XDFFA1/N1_XBOOTH/Xdffa1/M7_g N_VDD_XBOOTH/Xdffa1/M7_s
+ N_VDD_XBOOTH/Xdffa1/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXADDER/Xa000/Xao2/M36 N_XADDER/XA000/XAO2/N008_XADDER/Xa000/Xao2/M36_d
+ N_XADDER/XA000/OUT1_XADDER/Xa000/Xao2/M36_g
+ N_XADDER/XA000/XAO2/N007_XADDER/Xa000/Xao2/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXADDER/Xa01/Xrb1/M12 N_XADDER/XA01/XRB1/N003_XADDER/Xa01/Xrb1/M12_d
+ N_S[0]_XADDER/Xa01/Xrb1/M12_g N_VDD_XADDER/Xa01/Xrb1/M12_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/X_xor1/M5 N_XACCXOR/X_XOR1/N002_XACCXOR/X_xor1/M5_d
+ N_XACCXOR/DACC[1]_XACCXOR/X_xor1/M5_g
+ N_XACCXOR/X_XOR1/N001_XACCXOR/X_xor1/M5_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/X_xor2/M5 N_XACCXOR/X_XOR2/N002_XACCXOR/X_xor2/M5_d
+ N_XACCXOR/DACC[2]_XACCXOR/X_xor2/M5_g
+ N_XACCXOR/X_XOR2/N001_XACCXOR/X_xor2/M5_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/X_xor4/M5 N_XACCXOR/X_XOR4/N002_XACCXOR/X_xor4/M5_d
+ N_XACCXOR/DACC[4]_XACCXOR/X_xor4/M5_g
+ N_XACCXOR/X_XOR4/N001_XACCXOR/X_xor4/M5_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/X_xor6/M5 N_XACCXOR/X_XOR6/N002_XACCXOR/X_xor6/M5_d
+ N_XACCXOR/DACC[6]_XACCXOR/X_xor6/M5_g
+ N_XACCXOR/X_XOR6/N001_XACCXOR/X_xor6/M5_s N_VDD_XACCXOR/X_xor6/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/X_xor8/M5 N_XACCXOR/X_XOR8/N002_XACCXOR/X_xor8/M5_d
+ N_XACCXOR/DACC[8]_XACCXOR/X_xor8/M5_g
+ N_XACCXOR/X_XOR8/N001_XACCXOR/X_xor8/M5_s N_VDD_XACCXOR/X_xor6/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/X_xor10/M5 N_XACCXOR/X_XOR10/N002_XACCXOR/X_xor10/M5_d
+ N_XACCXOR/DACC[10]_XACCXOR/X_xor10/M5_g
+ N_XACCXOR/X_XOR10/N001_XACCXOR/X_xor10/M5_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa000/Xao2/M35 N_XADDER/XA000/XAO2/N007_XADDER/Xa000/Xao2/M35_d
+ N_XADDER/G0_XADDER/Xa000/Xao2/M35_g N_VDD_XADDER/Xa000/Xao2/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXADDER/Xa01/Xrb1/M11 N_XADDER/XA01/XRB1/N003_XADDER/Xa01/Xrb1/M11_d
+ N_GND_XADDER/Xa01/Xrb1/M11_g N_VDD_XADDER/Xa01/Xrb1/M11_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/X_xor1/M6 N_XACCXOR/X_XOR1/N001_XACCXOR/X_xor1/M6_d
+ N_DMODE_XACCXOR/X_xor1/M6_g N_VDD_XACCXOR/X_xor1/M6_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/X_xor2/M6 N_XACCXOR/X_XOR2/N001_XACCXOR/X_xor2/M6_d
+ N_DMODE_XACCXOR/X_xor2/M6_g N_VDD_XACCXOR/X_xor2/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/X_xor4/M6 N_XACCXOR/X_XOR4/N001_XACCXOR/X_xor4/M6_d
+ N_DMODE_XACCXOR/X_xor4/M6_g N_VDD_XACCXOR/X_xor4/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/X_xor6/M6 N_XACCXOR/X_XOR6/N001_XACCXOR/X_xor6/M6_d
+ N_DMODE_XACCXOR/X_xor6/M6_g N_VDD_XACCXOR/X_xor6/M6_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/X_xor8/M6 N_XACCXOR/X_XOR8/N001_XACCXOR/X_xor8/M6_d
+ N_DMODE_XACCXOR/X_xor8/M6_g N_VDD_XACCXOR/X_xor8/M6_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/X_xor10/M6 N_XACCXOR/X_XOR10/N001_XACCXOR/X_xor10/M6_d
+ N_DMODE_XACCXOR/X_xor10/M6_g N_VDD_XACCXOR/X_xor10/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mX02/xd21/M1 N_X02/XD21/P001_X02/xd21/M1_d N_OUT1[0]_X02/xd21/M1_g
+ N_VDD_X02/xd21/M1_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14
+ AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXADDER/Xa73/M4 N_OUT1[3]_XADDER/Xa73/M4_d N_XADDER/XA73/N002_XADDER/Xa73/M4_g
+ N_VDD_XADDER/Xa73/M4_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xdffa4/M10 N_XBOOTH/A_D[4]_XBOOTH/Xdffa4/M10_d
+ N_XBOOTH/XDFFA4/N3_XBOOTH/Xdffa4/M10_g N_VDD_XBOOTH/Xdffa4/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXBOOTH/Xdffa5/M10 N_A_D[5]_XBOOTH/Xdffa5/M10_d
+ N_XBOOTH/XDFFA5/N3_XBOOTH/Xdffa5/M10_g N_VDD_XBOOTH/Xdffa5/M10_s
+ N_VDD_XBOOTH/Xdffa5/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXBOOTH/Xdffa3/M10 N_A_D[3]_XBOOTH/Xdffa3/M10_d
+ N_XBOOTH/XDFFA3/N3_XBOOTH/Xdffa3/M10_g N_VDD_XBOOTH/Xdffa3/M10_s
+ N_VDD_XBOOTH/Xdffa5/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXBOOTH/Xdffa2/M10 N_XBOOTH/A_D[2]_XBOOTH/Xdffa2/M10_d
+ N_XBOOTH/XDFFA2/N3_XBOOTH/Xdffa2/M10_g N_VDD_XBOOTH/Xdffa2/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXBOOTH/Xdffa0/M10 N_XBOOTH/A_D[0]_XBOOTH/Xdffa0/M10_d
+ N_XBOOTH/XDFFA0/N3_XBOOTH/Xdffa0/M10_g N_VDD_XBOOTH/Xdffa0/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXBOOTH/Xdffa1/M10 N_A_D[1]_XBOOTH/Xdffa1/M10_d
+ N_XBOOTH/XDFFA1/N3_XBOOTH/Xdffa1/M10_g N_VDD_XBOOTH/Xdffa1/M10_s
+ N_VDD_XBOOTH/Xdffa1/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa000/Xao2/Xor1/M15 N_VDD_XADDER/Xa000/Xao2/Xor1/M15_d
+ N_XADDER/XA000/XAO2/N008_XADDER/Xa000/Xao2/Xor1/M15_g
+ N_XADDER/G00_XADDER/Xa000/Xao2/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mX02/xd21/M2 N_X02/XD21/N0_X02/xd21/M2_d N_CLK_X02/xd21/M2_g
+ N_X02/XD21/P001_X02/xd21/M2_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa01/Xrb1/Xand1/M15 N_VDD_XADDER/Xa01/Xrb1/Xand1/M15_d
+ N_XADDER/XA01/XRB1/N003_XADDER/Xa01/Xrb1/Xand1/M15_g
+ N_XADDER/G0_XADDER/Xa01/Xrb1/Xand1/M15_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXACCXOR/Xdffa12/M1 N_XACCXOR/XDFFA12/P001_XACCXOR/Xdffa12/M1_d
+ N_MODE_XACCXOR/Xdffa12/M1_g N_VDD_XACCXOR/Xdffa12/M1_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/Xdffa1/M10 N_XACCXOR/DACC[1]_XACCXOR/Xdffa1/M10_d
+ N_XACCXOR/XDFFA1/N3_XACCXOR/Xdffa1/M10_g N_VDD_XACCXOR/Xdffa1/M10_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/Xdffa2/M10 N_XACCXOR/DACC[2]_XACCXOR/Xdffa2/M10_d
+ N_XACCXOR/XDFFA2/N3_XACCXOR/Xdffa2/M10_g N_VDD_XACCXOR/Xdffa2/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/Xdffa4/M10 N_XACCXOR/DACC[4]_XACCXOR/Xdffa4/M10_d
+ N_XACCXOR/XDFFA4/N3_XACCXOR/Xdffa4/M10_g N_VDD_XACCXOR/Xdffa4/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/Xdffa6/M10 N_XACCXOR/DACC[6]_XACCXOR/Xdffa6/M10_d
+ N_XACCXOR/XDFFA6/N3_XACCXOR/Xdffa6/M10_g N_VDD_XACCXOR/Xdffa6/M10_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/Xdffa8/M10 N_XACCXOR/DACC[8]_XACCXOR/Xdffa8/M10_d
+ N_XACCXOR/XDFFA8/N3_XACCXOR/Xdffa8/M10_g N_VDD_XACCXOR/Xdffa8/M10_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/Xdffa10/M10 N_XACCXOR/DACC[10]_XACCXOR/Xdffa10/M10_d
+ N_XACCXOR/XDFFA10/N3_XACCXOR/Xdffa10/M10_g N_VDD_XACCXOR/Xdffa10/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa71/M6 N_XADDER/XA71/N001_XADDER/Xa71/M6_d
+ N_XADDER/G00_XADDER/Xa71/M6_g N_VDD_XADDER/Xa71/M6_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/Xdffa12/M2 N_XACCXOR/XDFFA12/N0_XACCXOR/Xdffa12/M2_d
+ N_CLK_XACCXOR/Xdffa12/M2_g N_XACCXOR/XDFFA12/P001_XACCXOR/Xdffa12/M2_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mX02/xd21/M4 N_X02/XD21/N1_X02/xd21/M4_d N_CLK_X02/xd21/M4_g N_VDD_X02/xd21/M4_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa71/M5 N_XADDER/XA71/N002_XADDER/Xa71/M5_d N_XADDER/P1_XADDER/Xa71/M5_g
+ N_XADDER/XA71/N001_XADDER/Xa71/M5_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=4.444e-13 AS=6.16e-14 PD=2.46e-06 PS=2.8e-07
mXADDER/Xa73/M5 N_XADDER/XA73/N002_XADDER/Xa73/M5_d N_XADDER/P3_XADDER/Xa73/M5_g
+ N_XADDER/XA73/N001_XADDER/Xa73/M5_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=4.444e-13 AS=6.16e-14 PD=2.46e-06 PS=2.8e-07
mXBOOTH/Xe2/M17 N_XBOOTH/XE2/_B_XBOOTH/Xe2/M17_d
+ N_XBOOTH/A_D[4]_XBOOTH/Xe2/M17_g N_VDD_XBOOTH/Xe2/M17_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe1/M17 N_XBOOTH/XE1/_B_XBOOTH/Xe1/M17_d
+ N_XBOOTH/A_D[2]_XBOOTH/Xe1/M17_g N_VDD_XBOOTH/Xe1/M17_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe0/M17 N_XBOOTH/XE0/_B_XBOOTH/Xe0/M17_d
+ N_XBOOTH/A_D[0]_XBOOTH/Xe0/M17_g N_VDD_XBOOTH/Xe0/M17_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa11/Xyb1/Xand1/M15 N_VDD_XADDER/Xa11/Xyb1/Xand1/M15_d
+ N_XADDER/XA11/XYB1/N003_XADDER/Xa11/Xyb1/Xand1/M15_g
+ N_XADDER/PP1_XADDER/Xa11/Xyb1/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa73/M6 N_XADDER/XA73/N001_XADDER/Xa73/M6_d
+ N_XADDER/GX6[0]_XADDER/Xa73/M6_g N_VDD_XADDER/Xa73/M6_s N_VDD_XADDER/Xa72/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXADDER/Xa02/Xrb2/M4 N_XADDER/P1_XADDER/Xa02/Xrb2/M4_d
+ N_XADDER/XA02/XRB2/N002_XADDER/Xa02/Xrb2/M4_g N_VDD_XADDER/Xa02/Xrb2/M4_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mX02/xd21/M7 N_X02/XD21/N3_X02/xd21/M7_d N_X02/XD21/N1_X02/xd21/M7_g
+ N_VDD_X02/xd21/M7_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa1/M7 N_XACCXOR/XDFFA1/N3_XACCXOR/Xdffa1/M7_d
+ N_XACCXOR/XDFFA1/N1_XACCXOR/Xdffa1/M7_g N_VDD_XACCXOR/Xdffa1/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa2/M7 N_XACCXOR/XDFFA2/N3_XACCXOR/Xdffa2/M7_d
+ N_XACCXOR/XDFFA2/N1_XACCXOR/Xdffa2/M7_g N_VDD_XACCXOR/Xdffa2/M7_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa4/M7 N_XACCXOR/XDFFA4/N3_XACCXOR/Xdffa4/M7_d
+ N_XACCXOR/XDFFA4/N1_XACCXOR/Xdffa4/M7_g N_VDD_XACCXOR/Xdffa4/M7_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa6/M7 N_XACCXOR/XDFFA6/N3_XACCXOR/Xdffa6/M7_d
+ N_XACCXOR/XDFFA6/N1_XACCXOR/Xdffa6/M7_g N_VDD_XACCXOR/Xdffa6/M7_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa8/M7 N_XACCXOR/XDFFA8/N3_XACCXOR/Xdffa8/M7_d
+ N_XACCXOR/XDFFA8/N1_XACCXOR/Xdffa8/M7_g N_VDD_XACCXOR/Xdffa8/M7_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa10/M7 N_XACCXOR/XDFFA10/N3_XACCXOR/Xdffa10/M7_d
+ N_XACCXOR/XDFFA10/N1_XACCXOR/Xdffa10/M7_g N_VDD_XACCXOR/Xdffa10/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe2/M16 N_XBOOTH/XE2/_A_XBOOTH/Xe2/M16_d N_A_D[5]_XBOOTH/Xe2/M16_g
+ N_VDD_XBOOTH/Xe2/M16_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.464e-13 AS=1.188e-13 PD=1.56e-06 PS=5.4e-07
mXBOOTH/Xe1/M16 N_XBOOTH/XE1/_A_XBOOTH/Xe1/M16_d N_A_D[3]_XBOOTH/Xe1/M16_g
+ N_VDD_XBOOTH/Xe1/M16_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.464e-13 AS=1.188e-13 PD=1.56e-06 PS=5.4e-07
mXBOOTH/Xe0/M16 N_XBOOTH/XE0/_A_XBOOTH/Xe0/M16_d N_A_D[1]_XBOOTH/Xe0/M16_g
+ N_VDD_XBOOTH/Xe0/M16_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.464e-13 AS=1.188e-13 PD=1.56e-06 PS=5.4e-07
mXACCXOR/Xdffa12/M4 N_XACCXOR/XDFFA12/N1_XACCXOR/Xdffa12/M4_d
+ N_CLK_XACCXOR/Xdffa12/M4_g N_VDD_XACCXOR/Xdffa12/M4_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa1/M4 N_XACCXOR/XDFFA1/N1_XACCXOR/Xdffa1/M4_d
+ N_CLK_XACCXOR/Xdffa1/M4_g N_VDD_XACCXOR/Xdffa1/M4_s N_VDD_XACCXOR/X_xor1/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa2/M4 N_XACCXOR/XDFFA2/N1_XACCXOR/Xdffa2/M4_d
+ N_CLK_XACCXOR/Xdffa2/M4_g N_VDD_XACCXOR/Xdffa2/M4_s N_VDD_XACCXOR/X_xor2/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa4/M4 N_XACCXOR/XDFFA4/N1_XACCXOR/Xdffa4/M4_d
+ N_CLK_XACCXOR/Xdffa4/M4_g N_VDD_XACCXOR/Xdffa4/M4_s N_VDD_XACCXOR/X_xor2/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa6/M4 N_XACCXOR/XDFFA6/N1_XACCXOR/Xdffa6/M4_d
+ N_CLK_XACCXOR/Xdffa6/M4_g N_VDD_XACCXOR/Xdffa6/M4_s N_VDD_XACCXOR/X_xor6/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa8/M4 N_XACCXOR/XDFFA8/N1_XACCXOR/Xdffa8/M4_d
+ N_CLK_XACCXOR/Xdffa8/M4_g N_VDD_XACCXOR/Xdffa8/M4_s N_VDD_XACCXOR/X_xor6/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa10/M4 N_XACCXOR/XDFFA10/N1_XACCXOR/Xdffa10/M4_d
+ N_CLK_XACCXOR/Xdffa10/M4_g N_VDD_XACCXOR/Xdffa10/M4_s N_VDD_XBOOTH/Xdffa4/M1_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa12/M7 N_XACCXOR/XDFFA12/N3_XACCXOR/Xdffa12/M7_d
+ N_XACCXOR/XDFFA12/N1_XACCXOR/Xdffa12/M7_g N_VDD_XACCXOR/Xdffa12/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa71/M4 N_OUT1[1]_XADDER/Xa71/M4_d N_XADDER/XA71/N002_XADDER/Xa71/M4_g
+ N_VDD_XADDER/Xa71/M4_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa11/Xyb1/M11 N_XADDER/XA11/XYB1/N003_XADDER/Xa11/Xyb1/M11_d
+ N_XADDER/P0_XADDER/Xa11/Xyb1/M11_g N_VDD_XADDER/Xa11/Xyb1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mX02/xd21/M10 N_OUT[0]_X02/xd21/M10_d N_X02/XD21/N3_X02/xd21/M10_g
+ N_VDD_X02/xd21/M10_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa02/Xrb2/M5 N_XADDER/XA02/XRB2/N001_XADDER/Xa02/Xrb2/M5_d
+ N_C[1]_XADDER/Xa02/Xrb2/M5_g N_VDD_XADDER/Xa02/Xrb2/M5_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.904e-13
+ PD=2.8e-07 PS=1.76e-06
mXBOOTH/Xe2/M10 N_noxref_1445_XBOOTH/Xe2/M10_d N_XBOOTH/XE2/_A_XBOOTH/Xe2/M10_g
+ N_VDD_XBOOTH/Xe2/M10_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe2/M13 N_XBOOTH/XE2/N002_XBOOTH/Xe2/M13_d N_A_D[5]_XBOOTH/Xe2/M13_g
+ N_noxref_1445_XBOOTH/Xe2/M13_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xe1/M13 N_XBOOTH/XE1/N002_XBOOTH/Xe1/M13_d N_A_D[3]_XBOOTH/Xe1/M13_g
+ N_noxref_1446_XBOOTH/Xe1/M13_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xe1/M10 N_noxref_1446_XBOOTH/Xe1/M10_d N_XBOOTH/XE1/_A_XBOOTH/Xe1/M10_g
+ N_VDD_XBOOTH/Xe1/M10_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe0/M10 N_noxref_1447_XBOOTH/Xe0/M10_d N_XBOOTH/XE0/_A_XBOOTH/Xe0/M10_g
+ N_VDD_XBOOTH/Xe0/M10_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe0/M13 N_XBOOTH/XE0/N002_XBOOTH/Xe0/M13_d N_A_D[1]_XBOOTH/Xe0/M13_g
+ N_noxref_1447_XBOOTH/Xe0/M13_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXADDER/Xa74/M4 N_OUT1[4]_XADDER/Xa74/M4_d N_XADDER/XA74/N002_XADDER/Xa74/M4_g
+ N_VDD_XADDER/Xa74/M4_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa11/Xyb1/M12 N_XADDER/XA11/XYB1/N003_XADDER/Xa11/Xyb1/M12_d
+ N_XADDER/P1_XADDER/Xa11/Xyb1/M12_g N_VDD_XADDER/Xa11/Xyb1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa02/Xrb2/M6 N_XADDER/XA02/XRB2/N002_XADDER/Xa02/Xrb2/M6_d
+ N_S[1]_XADDER/Xa02/Xrb2/M6_g N_XADDER/XA02/XRB2/N001_XADDER/Xa02/Xrb2/M6_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa1/M2 N_XACCXOR/XDFFA1/N0_XACCXOR/Xdffa1/M2_d
+ N_CLK_XACCXOR/Xdffa1/M2_g N_XACCXOR/XDFFA1/P001_XACCXOR/Xdffa1/M2_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa2/M2 N_XACCXOR/XDFFA2/N0_XACCXOR/Xdffa2/M2_d
+ N_CLK_XACCXOR/Xdffa2/M2_g N_XACCXOR/XDFFA2/P001_XACCXOR/Xdffa2/M2_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa4/M2 N_XACCXOR/XDFFA4/N0_XACCXOR/Xdffa4/M2_d
+ N_CLK_XACCXOR/Xdffa4/M2_g N_XACCXOR/XDFFA4/P001_XACCXOR/Xdffa4/M2_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa6/M2 N_XACCXOR/XDFFA6/N0_XACCXOR/Xdffa6/M2_d
+ N_CLK_XACCXOR/Xdffa6/M2_g N_XACCXOR/XDFFA6/P001_XACCXOR/Xdffa6/M2_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa8/M2 N_XACCXOR/XDFFA8/N0_XACCXOR/Xdffa8/M2_d
+ N_CLK_XACCXOR/Xdffa8/M2_g N_XACCXOR/XDFFA8/P001_XACCXOR/Xdffa8/M2_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa10/M2 N_XACCXOR/XDFFA10/N0_XACCXOR/Xdffa10/M2_d
+ N_CLK_XACCXOR/Xdffa10/M2_g N_XACCXOR/XDFFA10/P001_XACCXOR/Xdffa10/M2_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xe2/M11 N_noxref_1445_XBOOTH/Xe2/M11_d N_XBOOTH/A_D[4]_XBOOTH/Xe2/M11_g
+ N_VDD_XBOOTH/Xe2/M11_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=1.188e-13 PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xe2/M14 N_XBOOTH/XE2/N002_XBOOTH/Xe2/M14_d
+ N_XBOOTH/XE2/_B_XBOOTH/Xe2/M14_g N_noxref_1445_XBOOTH/Xe2/M14_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xe1/M14 N_XBOOTH/XE1/N002_XBOOTH/Xe1/M14_d
+ N_XBOOTH/XE1/_B_XBOOTH/Xe1/M14_g N_noxref_1446_XBOOTH/Xe1/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xe1/M11 N_noxref_1446_XBOOTH/Xe1/M11_d N_XBOOTH/A_D[2]_XBOOTH/Xe1/M11_g
+ N_VDD_XBOOTH/Xe1/M11_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=1.188e-13 PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xe0/M11 N_noxref_1447_XBOOTH/Xe0/M11_d N_XBOOTH/A_D[0]_XBOOTH/Xe0/M11_g
+ N_VDD_XBOOTH/Xe0/M11_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=1.188e-13 PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xe0/M14 N_XBOOTH/XE0/N002_XBOOTH/Xe0/M14_d
+ N_XBOOTH/XE0/_B_XBOOTH/Xe0/M14_g N_noxref_1447_XBOOTH/Xe0/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXACCXOR/Xdffa12/M10 N_DMODE_XACCXOR/Xdffa12/M10_d
+ N_XACCXOR/XDFFA12/N3_XACCXOR/Xdffa12/M10_g N_VDD_XACCXOR/Xdffa12/M10_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mX02/xd22/M1 N_X02/XD22/P001_X02/xd22/M1_d N_OUT1[1]_X02/xd22/M1_g
+ N_VDD_X02/xd22/M1_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14
+ AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXACCXOR/Xdffa1/M1 N_XACCXOR/XDFFA1/P001_XACCXOR/Xdffa1/M1_d
+ N_ACC[1]_XACCXOR/Xdffa1/M1_g N_VDD_XACCXOR/Xdffa1/M1_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/Xdffa2/M1 N_XACCXOR/XDFFA2/P001_XACCXOR/Xdffa2/M1_d
+ N_ACC[2]_XACCXOR/Xdffa2/M1_g N_VDD_XACCXOR/Xdffa2/M1_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/Xdffa4/M1 N_XACCXOR/XDFFA4/P001_XACCXOR/Xdffa4/M1_d
+ N_ACC[4]_XACCXOR/Xdffa4/M1_g N_VDD_XACCXOR/Xdffa4/M1_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/Xdffa6/M1 N_XACCXOR/XDFFA6/P001_XACCXOR/Xdffa6/M1_d
+ N_ACC[6]_XACCXOR/Xdffa6/M1_g N_VDD_XACCXOR/Xdffa6/M1_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/Xdffa8/M1 N_XACCXOR/XDFFA8/P001_XACCXOR/Xdffa8/M1_d
+ N_ACC[8]_XACCXOR/Xdffa8/M1_g N_VDD_XACCXOR/Xdffa8/M1_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/Xdffa10/M1 N_XACCXOR/XDFFA10/P001_XACCXOR/Xdffa10/M1_d
+ N_ACC[10]_XACCXOR/Xdffa10/M1_g N_VDD_XACCXOR/Xdffa10/M1_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXADDER/Xa62/Xao2/Xor1/M15 N_VDD_XADDER/Xa62/Xao2/Xor1/M15_d
+ N_XADDER/XA62/XAO2/N008_XADDER/Xa62/Xao2/Xor1/M15_g
+ N_XADDER/GX6[0]_XADDER/Xa62/Xao2/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mX02/xd22/M2 N_X02/XD22/N0_X02/xd22/M2_d N_CLK_X02/xd22/M2_g
+ N_X02/XD22/P001_X02/xd22/M2_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xe2/M12 N_noxref_1445_XBOOTH/Xe2/M12_d N_A_D[3]_XBOOTH/Xe2/M12_g
+ N_VDD_XBOOTH/Xe2/M12_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xe2/M15 N_XBOOTH/XE2/N002_XBOOTH/Xe2/M15_d
+ N_XBOOTH/XE2/_C_XBOOTH/Xe2/M15_g N_noxref_1445_XBOOTH/Xe2/M15_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe1/M15 N_XBOOTH/XE1/N002_XBOOTH/Xe1/M15_d
+ N_XBOOTH/XE1/_C_XBOOTH/Xe1/M15_g N_noxref_1446_XBOOTH/Xe1/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe1/M12 N_noxref_1446_XBOOTH/Xe1/M12_d N_A_D[1]_XBOOTH/Xe1/M12_g
+ N_VDD_XBOOTH/Xe1/M12_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xe0/M12 N_noxref_1447_XBOOTH/Xe0/M12_d N_GND_XBOOTH/Xe0/M12_g
+ N_VDD_XBOOTH/Xe0/M12_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=1.188e-13 AS=2.156e-13 PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xe0/M15 N_XBOOTH/XE0/N002_XBOOTH/Xe0/M15_d
+ N_XBOOTH/XE0/_C_XBOOTH/Xe0/M15_g N_noxref_1447_XBOOTH/Xe0/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa11/Xyb2/M12 N_XADDER/XA11/XYB2/N003_XADDER/Xa11/Xyb2/M12_d
+ N_XADDER/P1_XADDER/Xa11/Xyb2/M12_g N_VDD_XADDER/Xa11/Xyb2/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa02/Xrb1/M12 N_XADDER/XA02/XRB1/N003_XADDER/Xa02/Xrb1/M12_d
+ N_S[1]_XADDER/Xa02/Xrb1/M12_g N_VDD_XADDER/Xa02/Xrb1/M12_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa74/M5 N_XADDER/XA74/N002_XADDER/Xa74/M5_d N_XADDER/P4_XADDER/Xa74/M5_g
+ N_XADDER/XA74/N001_XADDER/Xa74/M5_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=4.444e-13 AS=6.16e-14 PD=2.46e-06 PS=2.8e-07
mXADDER/Xa62/Xao2/M35 N_XADDER/XA62/XAO2/N007_XADDER/Xa62/Xao2/M35_d
+ N_XADDER/G2_XADDER/Xa62/Xao2/M35_g N_VDD_XADDER/Xa62/Xao2/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXADDER/Xa11/Xyb2/M11 N_XADDER/XA11/XYB2/N003_XADDER/Xa11/Xyb2/M11_d
+ N_XADDER/G00_XADDER/Xa11/Xyb2/M11_g N_VDD_XADDER/Xa11/Xyb2/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mXACCXOR/Xdffa0/M1 N_XACCXOR/XDFFA0/P001_XACCXOR/Xdffa0/M1_d
+ N_ACC[0]_XACCXOR/Xdffa0/M1_g N_VDD_XACCXOR/Xdffa0/M1_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/Xdffa3/M1 N_XACCXOR/XDFFA3/P001_XACCXOR/Xdffa3/M1_d
+ N_ACC[3]_XACCXOR/Xdffa3/M1_g N_VDD_XACCXOR/Xdffa3/M1_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/Xdffa5/M1 N_XACCXOR/XDFFA5/P001_XACCXOR/Xdffa5/M1_d
+ N_ACC[5]_XACCXOR/Xdffa5/M1_g N_VDD_XACCXOR/Xdffa5/M1_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/Xdffa7/M1 N_XACCXOR/XDFFA7/P001_XACCXOR/Xdffa7/M1_d
+ N_ACC[7]_XACCXOR/Xdffa7/M1_g N_VDD_XACCXOR/Xdffa7/M1_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/Xdffa9/M1 N_XACCXOR/XDFFA9/P001_XACCXOR/Xdffa9/M1_d
+ N_ACC[9]_XACCXOR/Xdffa9/M1_g N_VDD_XACCXOR/Xdffa9/M1_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/Xdffa11/M1 N_XACCXOR/XDFFA11/P001_XACCXOR/Xdffa11/M1_d
+ N_ACC[11]_XACCXOR/Xdffa11/M1_g N_VDD_XACCXOR/Xdffa11/M1_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXADDER/Xa74/M6 N_XADDER/XA74/N001_XADDER/Xa74/M6_d
+ N_XADDER/GGG3_XADDER/Xa74/M6_g N_VDD_XADDER/Xa74/M6_s N_VDD_XADDER/Xa72/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXADDER/Xa02/Xrb1/M11 N_XADDER/XA02/XRB1/N003_XADDER/Xa02/Xrb1/M11_d
+ N_C[1]_XADDER/Xa02/Xrb1/M11_g N_VDD_XADDER/Xa02/Xrb1/M11_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd22/M4 N_X02/XD22/N1_X02/xd22/M4_d N_CLK_X02/xd22/M4_g N_VDD_X02/xd22/M4_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa62/Xao2/M36 N_XADDER/XA62/XAO2/N008_XADDER/Xa62/Xao2/M36_d
+ N_XADDER/XA62/OUT1_XADDER/Xa62/Xao2/M36_g
+ N_XADDER/XA62/XAO2/N007_XADDER/Xa62/Xao2/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXBOOTH/Xe2/M18 N_XBOOTH/XE2/_C_XBOOTH/Xe2/M18_d N_A_D[3]_XBOOTH/Xe2/M18_g
+ N_VDD_XBOOTH/Xe2/M18_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.41576e-13 PD=1.42e-06 PS=5.69412e-07
mXBOOTH/Xe1/M18 N_XBOOTH/XE1/_C_XBOOTH/Xe1/M18_d N_A_D[1]_XBOOTH/Xe1/M18_g
+ N_VDD_XBOOTH/Xe1/M18_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.41576e-13 PD=1.42e-06 PS=5.69412e-07
mXBOOTH/Xe0/M18 N_XBOOTH/XE0/_C_XBOOTH/Xe0/M18_d N_GND_XBOOTH/Xe0/M18_g
+ N_VDD_XBOOTH/Xe0/M18_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.41576e-13 PD=1.42e-06 PS=5.69412e-07
mXACCXOR/Xdffa0/M2 N_XACCXOR/XDFFA0/N0_XACCXOR/Xdffa0/M2_d
+ N_CLK_XACCXOR/Xdffa0/M2_g N_XACCXOR/XDFFA0/P001_XACCXOR/Xdffa0/M2_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa3/M2 N_XACCXOR/XDFFA3/N0_XACCXOR/Xdffa3/M2_d
+ N_CLK_XACCXOR/Xdffa3/M2_g N_XACCXOR/XDFFA3/P001_XACCXOR/Xdffa3/M2_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa5/M2 N_XACCXOR/XDFFA5/N0_XACCXOR/Xdffa5/M2_d
+ N_CLK_XACCXOR/Xdffa5/M2_g N_XACCXOR/XDFFA5/P001_XACCXOR/Xdffa5/M2_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa7/M2 N_XACCXOR/XDFFA7/N0_XACCXOR/Xdffa7/M2_d
+ N_CLK_XACCXOR/Xdffa7/M2_g N_XACCXOR/XDFFA7/P001_XACCXOR/Xdffa7/M2_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa9/M2 N_XACCXOR/XDFFA9/N0_XACCXOR/Xdffa9/M2_d
+ N_CLK_XACCXOR/Xdffa9/M2_g N_XACCXOR/XDFFA9/P001_XACCXOR/Xdffa9/M2_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXACCXOR/Xdffa11/M2 N_XACCXOR/XDFFA11/N0_XACCXOR/Xdffa11/M2_d
+ N_CLK_XACCXOR/Xdffa11/M2_g N_XACCXOR/XDFFA11/P001_XACCXOR/Xdffa11/M2_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mX02/xd22/M7 N_X02/XD22/N3_X02/xd22/M7_d N_X02/XD22/N1_X02/xd22/M7_g
+ N_VDD_X02/xd22/M7_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe2/M20 N_XBOOTH/D2_XBOOTH/Xe2/M20_d N_XBOOTH/XE2/N002_XBOOTH/Xe2/M20_g
+ N_VDD_XBOOTH/Xe2/M20_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.8e-07
+ AD=2.842e-13 AS=1.86624e-13 PD=1.56e-06 PS=7.50588e-07
mXBOOTH/Xe1/M20 N_XBOOTH/D1_XBOOTH/Xe1/M20_d N_XBOOTH/XE1/N002_XBOOTH/Xe1/M20_g
+ N_VDD_XBOOTH/Xe1/M20_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=5.8e-07
+ AD=2.842e-13 AS=1.86624e-13 PD=1.56e-06 PS=7.50588e-07
mXBOOTH/Xe0/M20 N_XBOOTH/D0_XBOOTH/Xe0/M20_d N_XBOOTH/XE0/N002_XBOOTH/Xe0/M20_g
+ N_VDD_XBOOTH/Xe0/M20_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=5.8e-07
+ AD=2.842e-13 AS=1.86624e-13 PD=1.56e-06 PS=7.50588e-07
mXADDER/Xa11/Xyb2/Xand1/M15 N_VDD_XADDER/Xa11/Xyb2/Xand1/M15_d
+ N_XADDER/XA11/XYB2/N003_XADDER/Xa11/Xyb2/Xand1/M15_g
+ N_XADDER/XA11/T1_XADDER/Xa11/Xyb2/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa02/Xrb1/Xand1/M15 N_VDD_XADDER/Xa02/Xrb1/Xand1/M15_d
+ N_XADDER/XA02/XRB1/N003_XADDER/Xa02/Xrb1/Xand1/M15_g
+ N_XADDER/G1_XADDER/Xa02/Xrb1/Xand1/M15_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa62/Xao1/Xand1/M15 N_VDD_XADDER/Xa62/Xao1/Xand1/M15_d
+ N_XADDER/XA62/XAO1/N003_XADDER/Xa62/Xao1/Xand1/M15_g
+ N_XADDER/XA62/OUT1_XADDER/Xa62/Xao1/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXACCXOR/Xdffa0/M4 N_XACCXOR/XDFFA0/N1_XACCXOR/Xdffa0/M4_d
+ N_CLK_XACCXOR/Xdffa0/M4_g N_VDD_XACCXOR/Xdffa0/M4_s N_VDD_XACCXOR/X_xor1/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa3/M4 N_XACCXOR/XDFFA3/N1_XACCXOR/Xdffa3/M4_d
+ N_CLK_XACCXOR/Xdffa3/M4_g N_VDD_XACCXOR/Xdffa3/M4_s N_VDD_XACCXOR/X_xor2/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa5/M4 N_XACCXOR/XDFFA5/N1_XACCXOR/Xdffa5/M4_d
+ N_CLK_XACCXOR/Xdffa5/M4_g N_VDD_XACCXOR/Xdffa5/M4_s N_VDD_XACCXOR/X_xor2/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa7/M4 N_XACCXOR/XDFFA7/N1_XACCXOR/Xdffa7/M4_d
+ N_CLK_XACCXOR/Xdffa7/M4_g N_VDD_XACCXOR/Xdffa7/M4_s N_VDD_XACCXOR/X_xor6/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa9/M4 N_XACCXOR/XDFFA9/N1_XACCXOR/Xdffa9/M4_d
+ N_CLK_XACCXOR/Xdffa9/M4_g N_VDD_XACCXOR/Xdffa9/M4_s N_VDD_XACCXOR/X_xor6/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa11/M4 N_XACCXOR/XDFFA11/N1_XACCXOR/Xdffa11/M4_d
+ N_CLK_XACCXOR/Xdffa11/M4_g N_VDD_XACCXOR/Xdffa11/M4_s N_VDD_XBOOTH/Xdffa4/M1_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mX02/xd22/M10 N_OUT[1]_X02/xd22/M10_d N_X02/XD22/N3_X02/xd22/M10_g
+ N_VDD_X02/xd22/M10_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXACCXOR/Xdffa0/M7 N_XACCXOR/XDFFA0/N3_XACCXOR/Xdffa0/M7_d
+ N_XACCXOR/XDFFA0/N1_XACCXOR/Xdffa0/M7_g N_VDD_XACCXOR/Xdffa0/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa3/M7 N_XACCXOR/XDFFA3/N3_XACCXOR/Xdffa3/M7_d
+ N_XACCXOR/XDFFA3/N1_XACCXOR/Xdffa3/M7_g N_VDD_XACCXOR/Xdffa3/M7_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa5/M7 N_XACCXOR/XDFFA5/N3_XACCXOR/Xdffa5/M7_d
+ N_XACCXOR/XDFFA5/N1_XACCXOR/Xdffa5/M7_g N_VDD_XACCXOR/Xdffa5/M7_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa7/M7 N_XACCXOR/XDFFA7/N3_XACCXOR/Xdffa7/M7_d
+ N_XACCXOR/XDFFA7/N1_XACCXOR/Xdffa7/M7_g N_VDD_XACCXOR/Xdffa7/M7_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa9/M7 N_XACCXOR/XDFFA9/N3_XACCXOR/Xdffa9/M7_d
+ N_XACCXOR/XDFFA9/N1_XACCXOR/Xdffa9/M7_g N_VDD_XACCXOR/Xdffa9/M7_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/Xdffa11/M7 N_XACCXOR/XDFFA11/N3_XACCXOR/Xdffa11/M7_d
+ N_XACCXOR/XDFFA11/N1_XACCXOR/Xdffa11/M7_g N_VDD_XACCXOR/Xdffa11/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xe2/M26 N_XBOOTH/XE2/N003_XBOOTH/Xe2/M26_d N_A_D[3]_XBOOTH/Xe2/M26_g
+ N_VDD_XBOOTH/Xe2/M26_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xe1/M26 N_XBOOTH/XE1/N003_XBOOTH/Xe1/M26_d N_A_D[1]_XBOOTH/Xe1/M26_g
+ N_VDD_XBOOTH/Xe1/M26_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xe0/M26 N_XBOOTH/XE0/N003_XBOOTH/Xe0/M26_d N_GND_XBOOTH/Xe0/M26_g
+ N_VDD_XBOOTH/Xe0/M26_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXADDER/Xa11/Xyb3/M36 N_XADDER/XA11/XYB3/N008_XADDER/Xa11/Xyb3/M36_d
+ N_XADDER/XA11/T1_XADDER/Xa11/Xyb3/M36_g
+ N_XADDER/XA11/XYB3/N007_XADDER/Xa11/Xyb3/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXADDER/Xa03/Xrb2/M4 N_XADDER/P2_XADDER/Xa03/Xrb2/M4_d
+ N_XADDER/XA03/XRB2/N002_XADDER/Xa03/Xrb2/M4_g N_VDD_XADDER/Xa03/Xrb2/M4_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xe2/M25 N_XBOOTH/XE2/N004_XBOOTH/Xe2/M25_d
+ N_XBOOTH/A_D[4]_XBOOTH/Xe2/M25_g N_XBOOTH/XE2/N003_XBOOTH/Xe2/M25_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xe1/M25 N_XBOOTH/XE1/N004_XBOOTH/Xe1/M25_d
+ N_XBOOTH/A_D[2]_XBOOTH/Xe1/M25_g N_XBOOTH/XE1/N003_XBOOTH/Xe1/M25_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xe0/M25 N_XBOOTH/XE0/N004_XBOOTH/Xe0/M25_d
+ N_XBOOTH/A_D[0]_XBOOTH/Xe0/M25_g N_XBOOTH/XE0/N003_XBOOTH/Xe0/M25_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa62/Xao1/M12 N_XADDER/XA62/XAO1/N003_XADDER/Xa62/Xao1/M12_d
+ N_XADDER/P2_XADDER/Xa62/Xao1/M12_g N_VDD_XADDER/Xa62/Xao1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.288e-13 AS=1.474e-13
+ PD=1.48e-06 PS=6.7e-07
mXADDER/Xa11/Xyb3/M35 N_XADDER/XA11/XYB3/N007_XADDER/Xa11/Xyb3/M35_d
+ N_XADDER/G1_XADDER/Xa11/Xyb3/M35_g N_VDD_XADDER/Xa11/Xyb3/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mX02/xd23/M1 N_X02/XD23/P001_X02/xd23/M1_d N_OUT1[2]_X02/xd23/M1_g
+ N_VDD_X02/xd23/M1_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14
+ AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXACCXOR/Xdffa0/M10 N_XACCXOR/DACC[0]_XACCXOR/Xdffa0/M10_d
+ N_XACCXOR/XDFFA0/N3_XACCXOR/Xdffa0/M10_g N_VDD_XACCXOR/Xdffa0/M10_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/Xdffa3/M10 N_XACCXOR/DACC[3]_XACCXOR/Xdffa3/M10_d
+ N_XACCXOR/XDFFA3/N3_XACCXOR/Xdffa3/M10_g N_VDD_XACCXOR/Xdffa3/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/Xdffa5/M10 N_XACCXOR/DACC[5]_XACCXOR/Xdffa5/M10_d
+ N_XACCXOR/XDFFA5/N3_XACCXOR/Xdffa5/M10_g N_VDD_XACCXOR/Xdffa5/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/Xdffa7/M10 N_XACCXOR/DACC[7]_XACCXOR/Xdffa7/M10_d
+ N_XACCXOR/XDFFA7/N3_XACCXOR/Xdffa7/M10_g N_VDD_XACCXOR/Xdffa7/M10_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/Xdffa9/M10 N_XACCXOR/DACC[9]_XACCXOR/Xdffa9/M10_d
+ N_XACCXOR/XDFFA9/N3_XACCXOR/Xdffa9/M10_g N_VDD_XACCXOR/Xdffa9/M10_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/Xdffa11/M10 N_XACCXOR/DACC[11]_XACCXOR/Xdffa11/M10_d
+ N_XACCXOR/XDFFA11/N3_XACCXOR/Xdffa11/M10_g N_VDD_XACCXOR/Xdffa11/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa62/Xao1/M11 N_XADDER/XA62/XAO1/N003_XADDER/Xa62/Xao1/M11_d
+ N_XADDER/GG1_XADDER/Xa62/Xao1/M11_g N_VDD_XADDER/Xa62/Xao1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.474e-13
+ PD=1.42e-06 PS=6.7e-07
mXADDER/Xa11/Xyb3/Xor1/M15 N_VDD_XADDER/Xa11/Xyb3/Xor1/M15_d
+ N_XADDER/XA11/XYB3/N008_XADDER/Xa11/Xyb3/Xor1/M15_g
+ N_XADDER/GG1_XADDER/Xa11/Xyb3/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mX02/xd23/M2 N_X02/XD23/N0_X02/xd23/M2_d N_CLK_X02/xd23/M2_g
+ N_X02/XD23/P001_X02/xd23/M2_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa03/Xrb2/M5 N_XADDER/XA03/XRB2/N001_XADDER/Xa03/Xrb2/M5_d
+ N_C[2]_XADDER/Xa03/Xrb2/M5_g N_VDD_XADDER/Xa03/Xrb2/M5_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.904e-13
+ PD=2.8e-07 PS=1.76e-06
mXCSA/Xdffmod/M1 N_XCSA/XDFFMOD/P001_XCSA/Xdffmod/M1_d N_DMODE_XCSA/Xdffmod/M1_g
+ N_VDD_XCSA/Xdffmod/M1_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa12/M1 N_XCSA/XDFFA12/P001_XCSA/Xdffa12/M1_d
+ N_XCSA/LV3_S[0]_XCSA/Xdffa12/M1_g N_VDD_XCSA/Xdffa12/M1_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xe2/M24 N_XBOOTH/S2_XBOOTH/Xe2/M24_d N_XBOOTH/XE2/N004_XBOOTH/Xe2/M24_g
+ N_VDD_XBOOTH/Xe2/M24_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.8e-07
+ AD=2.842e-13 AS=2.842e-13 PD=1.56e-06 PS=1.56e-06
mXBOOTH/Xe1/M24 N_XBOOTH/S1_XBOOTH/Xe1/M24_d N_XBOOTH/XE1/N004_XBOOTH/Xe1/M24_g
+ N_VDD_XBOOTH/Xe1/M24_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=5.8e-07
+ AD=2.842e-13 AS=2.842e-13 PD=1.56e-06 PS=1.56e-06
mXBOOTH/Xe0/M24 N_XBOOTH/S0_XBOOTH/Xe0/M24_d N_XBOOTH/XE0/N004_XBOOTH/Xe0/M24_g
+ N_VDD_XBOOTH/Xe0/M24_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=5.8e-07
+ AD=2.842e-13 AS=2.842e-13 PD=1.56e-06 PS=1.56e-06
mXADDER/Xa03/Xrb2/M6 N_XADDER/XA03/XRB2/N002_XADDER/Xa03/Xrb2/M6_d
+ N_S[2]_XADDER/Xa03/Xrb2/M6_g N_XADDER/XA03/XRB2/N001_XADDER/Xa03/Xrb2/M6_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffmod/M2 N_XCSA/XDFFMOD/N0_XCSA/Xdffmod/M2_d N_CLK_XCSA/Xdffmod/M2_g
+ N_XCSA/XDFFMOD/P001_XCSA/Xdffmod/M2_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa12/M2 N_XCSA/XDFFA12/N0_XCSA/Xdffa12/M2_d N_CLK_XCSA/Xdffa12/M2_g
+ N_XCSA/XDFFA12/P001_XCSA/Xdffa12/M2_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa23/Xao1/M11 N_XADDER/XA23/XAO1/N003_XADDER/Xa23/Xao1/M11_d
+ N_XADDER/GG1_XADDER/Xa23/Xao1/M11_g N_VDD_XADDER/Xa23/Xao1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.474e-13
+ PD=1.42e-06 PS=6.7e-07
mXACCXOR/X_xor0/M6 N_XACCXOR/X_XOR0/N001_XACCXOR/X_xor0/M6_d
+ N_DMODE_XACCXOR/X_xor0/M6_g N_VDD_XACCXOR/X_xor0/M6_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/X_xor3/M6 N_XACCXOR/X_XOR3/N001_XACCXOR/X_xor3/M6_d
+ N_DMODE_XACCXOR/X_xor3/M6_g N_VDD_XACCXOR/X_xor3/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/X_xor5/M6 N_XACCXOR/X_XOR5/N001_XACCXOR/X_xor5/M6_d
+ N_DMODE_XACCXOR/X_xor5/M6_g N_VDD_XACCXOR/X_xor5/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/X_xor7/M6 N_XACCXOR/X_XOR7/N001_XACCXOR/X_xor7/M6_d
+ N_DMODE_XACCXOR/X_xor7/M6_g N_VDD_XACCXOR/X_xor7/M6_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/X_xor9/M6 N_XACCXOR/X_XOR9/N001_XACCXOR/X_xor9/M6_d
+ N_DMODE_XACCXOR/X_xor9/M6_g N_VDD_XACCXOR/X_xor9/M6_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXACCXOR/X_xor11/M6 N_XACCXOR/X_XOR11/N001_XACCXOR/X_xor11/M6_d
+ N_DMODE_XACCXOR/X_xor11/M6_g N_VDD_XACCXOR/X_xor11/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mX02/xd23/M4 N_X02/XD23/N1_X02/xd23/M4_d N_CLK_X02/xd23/M4_g N_VDD_X02/xd23/M4_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXACCXOR/X_xor0/M5 N_XACCXOR/X_XOR0/N002_XACCXOR/X_xor0/M5_d
+ N_XACCXOR/DACC[0]_XACCXOR/X_xor0/M5_g
+ N_XACCXOR/X_XOR0/N001_XACCXOR/X_xor0/M5_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/X_xor3/M5 N_XACCXOR/X_XOR3/N002_XACCXOR/X_xor3/M5_d
+ N_XACCXOR/DACC[3]_XACCXOR/X_xor3/M5_g
+ N_XACCXOR/X_XOR3/N001_XACCXOR/X_xor3/M5_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/X_xor5/M5 N_XACCXOR/X_XOR5/N002_XACCXOR/X_xor5/M5_d
+ N_XACCXOR/DACC[5]_XACCXOR/X_xor5/M5_g
+ N_XACCXOR/X_XOR5/N001_XACCXOR/X_xor5/M5_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/X_xor7/M5 N_XACCXOR/X_XOR7/N002_XACCXOR/X_xor7/M5_d
+ N_XACCXOR/DACC[7]_XACCXOR/X_xor7/M5_g
+ N_XACCXOR/X_XOR7/N001_XACCXOR/X_xor7/M5_s N_VDD_XACCXOR/X_xor6/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/X_xor9/M5 N_XACCXOR/X_XOR9/N002_XACCXOR/X_xor9/M5_d
+ N_XACCXOR/DACC[9]_XACCXOR/X_xor9/M5_g
+ N_XACCXOR/X_XOR9/N001_XACCXOR/X_xor9/M5_s N_VDD_XACCXOR/X_xor6/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXACCXOR/X_xor11/M5 N_XACCXOR/X_XOR11/N002_XACCXOR/X_xor11/M5_d
+ N_XACCXOR/DACC[11]_XACCXOR/X_xor11/M5_g
+ N_XACCXOR/X_XOR11/N001_XACCXOR/X_xor11/M5_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa13/Xyb1/Xand1/M15 N_VDD_XADDER/Xa13/Xyb1/Xand1/M15_d
+ N_XADDER/XA13/XYB1/N003_XADDER/Xa13/Xyb1/Xand1/M15_g
+ N_XADDER/PP3_XADDER/Xa13/Xyb1/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa23/Xao1/M12 N_XADDER/XA23/XAO1/N003_XADDER/Xa23/Xao1/M12_d
+ N_XADDER/PP3_XADDER/Xa23/Xao1/M12_g N_VDD_XADDER/Xa23/Xao1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.288e-13 AS=1.474e-13
+ PD=1.48e-06 PS=6.7e-07
mXCSA/Xdffmod/M4 N_XCSA/XDFFMOD/N1_XCSA/Xdffmod/M4_d N_CLK_XCSA/Xdffmod/M4_g
+ N_VDD_XCSA/Xdffmod/M4_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa12/M4 N_XCSA/XDFFA12/N1_XCSA/Xdffa12/M4_d N_CLK_XCSA/Xdffa12/M4_g
+ N_VDD_XCSA/Xdffa12/M4_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mX02/xd23/M7 N_X02/XD23/N3_X02/xd23/M7_d N_X02/XD23/N1_X02/xd23/M7_g
+ N_VDD_X02/xd23/M7_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXADDER/Xa03/Xrb1/M12 N_XADDER/XA03/XRB1/N003_XADDER/Xa03/Xrb1/M12_d
+ N_S[2]_XADDER/Xa03/Xrb1/M12_g N_VDD_XADDER/Xa03/Xrb1/M12_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel20/M8 N_XBOOTH/XSEL20/N002_XBOOTH/Xsel20/M8_d
+ N_GND_XBOOTH/Xsel20/M8_g N_noxref_1508_XBOOTH/Xsel20/M8_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel10/M8 N_XBOOTH/XSEL10/N002_XBOOTH/Xsel10/M8_d
+ N_GND_XBOOTH/Xsel10/M8_g N_noxref_1509_XBOOTH/Xsel10/M8_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel00/M8 N_XBOOTH/XSEL00/N002_XBOOTH/Xsel00/M8_d
+ N_GND_XBOOTH/Xsel00/M8_g N_noxref_1510_XBOOTH/Xsel00/M8_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/Xdffmod/M7 N_XCSA/XDFFMOD/N3_XCSA/Xdffmod/M7_d
+ N_XCSA/XDFFMOD/N1_XCSA/Xdffmod/M7_g N_VDD_XCSA/Xdffmod/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa12/M7 N_XCSA/XDFFA12/N3_XCSA/Xdffa12/M7_d
+ N_XCSA/XDFFA12/N1_XCSA/Xdffa12/M7_g N_VDD_XCSA/Xdffa12/M7_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa03/Xrb1/M11 N_XADDER/XA03/XRB1/N003_XADDER/Xa03/Xrb1/M11_d
+ N_C[2]_XADDER/Xa03/Xrb1/M11_g N_VDD_XADDER/Xa03/Xrb1/M11_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel20/M6 N_XBOOTH/XSEL20/N002_XBOOTH/Xsel20/M6_d
+ N_XBOOTH/D2_XBOOTH/Xsel20/M6_g N_noxref_1508_XBOOTH/Xsel20/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel10/M6 N_XBOOTH/XSEL10/N002_XBOOTH/Xsel10/M6_d
+ N_XBOOTH/D1_XBOOTH/Xsel10/M6_g N_noxref_1509_XBOOTH/Xsel10/M6_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel00/M6 N_XBOOTH/XSEL00/N002_XBOOTH/Xsel00/M6_d
+ N_XBOOTH/D0_XBOOTH/Xsel00/M6_g N_noxref_1510_XBOOTH/Xsel00/M6_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXADDER/Xa13/Xyb1/M11 N_XADDER/XA13/XYB1/N003_XADDER/Xa13/Xyb1/M11_d
+ N_XADDER/P2_XADDER/Xa13/Xyb1/M11_g N_VDD_XADDER/Xa13/Xyb1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mXACCXOR/X_xor0/M4 N_CACC[0]_XACCXOR/X_xor0/M4_d
+ N_XACCXOR/X_XOR0/N002_XACCXOR/X_xor0/M4_g N_VDD_XACCXOR/X_xor0/M4_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor3/M4 N_CACC[3]_XACCXOR/X_xor3/M4_d
+ N_XACCXOR/X_XOR3/N002_XACCXOR/X_xor3/M4_g N_VDD_XACCXOR/X_xor3/M4_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor5/M4 N_CACC[5]_XACCXOR/X_xor5/M4_d
+ N_XACCXOR/X_XOR5/N002_XACCXOR/X_xor5/M4_g N_VDD_XACCXOR/X_xor5/M4_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor7/M4 N_CACC[7]_XACCXOR/X_xor7/M4_d
+ N_XACCXOR/X_XOR7/N002_XACCXOR/X_xor7/M4_g N_VDD_XACCXOR/X_xor7/M4_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor9/M4 N_CACC[9]_XACCXOR/X_xor9/M4_d
+ N_XACCXOR/X_XOR9/N002_XACCXOR/X_xor9/M4_g N_VDD_XACCXOR/X_xor9/M4_s
+ N_VDD_XACCXOR/X_xor6/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXACCXOR/X_xor11/M4 N_CACC[11]_XACCXOR/X_xor11/M4_d
+ N_XACCXOR/X_XOR11/N002_XACCXOR/X_xor11/M4_g N_VDD_XACCXOR/X_xor11/M4_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa23/Xao1/Xand1/M15 N_VDD_XADDER/Xa23/Xao1/Xand1/M15_d
+ N_XADDER/XA23/XAO1/N003_XADDER/Xa23/Xao1/Xand1/M15_g
+ N_XADDER/XA23/OUT1_XADDER/Xa23/Xao1/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd23/M10 N_OUT[2]_X02/xd23/M10_d N_X02/XD23/N3_X02/xd23/M10_g
+ N_VDD_X02/xd23/M10_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel20/M7 N_noxref_1508_XBOOTH/Xsel20/M7_d
+ N_XBOOTH/S2_XBOOTH/Xsel20/M7_g N_VDD_XBOOTH/Xsel20/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel10/M7 N_noxref_1509_XBOOTH/Xsel10/M7_d
+ N_XBOOTH/S1_XBOOTH/Xsel10/M7_g N_VDD_XBOOTH/Xsel10/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel00/M7 N_noxref_1510_XBOOTH/Xsel00/M7_d
+ N_XBOOTH/S0_XBOOTH/Xsel00/M7_g N_VDD_XBOOTH/Xsel00/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXADDER/Xa13/Xyb1/M12 N_XADDER/XA13/XYB1/N003_XADDER/Xa13/Xyb1/M12_d
+ N_XADDER/P3_XADDER/Xa13/Xyb1/M12_g N_VDD_XADDER/Xa13/Xyb1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffmod/M10 N_CIN_XCSA/Xdffmod/M10_d N_XCSA/XDFFMOD/N3_XCSA/Xdffmod/M10_g
+ N_VDD_XCSA/Xdffmod/M10_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa12/M10 N_S[0]_XCSA/Xdffa12/M10_d N_XCSA/XDFFA12/N3_XCSA/Xdffa12/M10_g
+ N_VDD_XCSA/Xdffa12/M10_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa03/Xrb1/Xand1/M15 N_VDD_XADDER/Xa03/Xrb1/Xand1/M15_d
+ N_XADDER/XA03/XRB1/N003_XADDER/Xa03/Xrb1/Xand1/M15_g
+ N_XADDER/G2_XADDER/Xa03/Xrb1/Xand1/M15_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel20/M9 N_noxref_1508_XBOOTH/Xsel20/M9_d
+ N_XBOOTH/B_D[0]_XBOOTH/Xsel20/M9_g N_VDD_XBOOTH/Xsel20/M9_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel10/M9 N_noxref_1509_XBOOTH/Xsel10/M9_d
+ N_XBOOTH/B_D[0]_XBOOTH/Xsel10/M9_g N_VDD_XBOOTH/Xsel10/M9_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel00/M9 N_noxref_1510_XBOOTH/Xsel00/M9_d
+ N_XBOOTH/B_D[0]_XBOOTH/Xsel00/M9_g N_VDD_XBOOTH/Xsel00/M9_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xdffb0/M1 N_XBOOTH/XDFFB0/P001_XBOOTH/Xdffb0/M1_d
+ N_B[0]_XBOOTH/Xdffb0/M1_g N_VDD_XBOOTH/Xdffb0/M1_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=7.7e-14 AS=2.695e-13 PD=2.8e-07 PS=1.53e-06
mXADDER/Xa23/Xao2/M36 N_XADDER/XA23/XAO2/N008_XADDER/Xa23/Xao2/M36_d
+ N_XADDER/XA23/OUT1_XADDER/Xa23/Xao2/M36_g
+ N_XADDER/XA23/XAO2/N007_XADDER/Xa23/Xao2/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mX02/xd24/M1 N_X02/XD24/P001_X02/xd24/M1_d N_OUT1[3]_X02/xd24/M1_g
+ N_VDD_X02/xd24/M1_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14
+ AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xdffb0/M2 N_XBOOTH/XDFFB0/N0_XBOOTH/Xdffb0/M2_d N_CLK_XBOOTH/Xdffb0/M2_g
+ N_XBOOTH/XDFFB0/P001_XBOOTH/Xdffb0/M2_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=7.7e-14 PD=1.53e-06 PS=2.8e-07
mXCSA/X_LV1_HA0/X_xor/M4 N_XCSA/LV1_S[2]_XCSA/X_LV1_HA0/X_xor/M4_d
+ N_XCSA/X_LV1_HA0/X_XOR/N002_XCSA/X_LV1_HA0/X_xor/M4_g
+ N_VDD_XCSA/X_LV1_HA0/X_xor/M4_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_HA0/M13 N_XCSA/LV1_C[3]_XCSA/X_LV1_HA0/M13_d
+ N_XCSA/X_LV1_HA0/N001_XCSA/X_LV1_HA0/M13_g N_VDD_XCSA/X_LV1_HA0/M13_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mX02/xd24/M2 N_X02/XD24/N0_X02/xd24/M2_d N_CLK_X02/xd24/M2_g
+ N_X02/XD24/P001_X02/xd24/M2_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa13/Xyb2/M12 N_XADDER/XA13/XYB2/N003_XADDER/Xa13/Xyb2/M12_d
+ N_XADDER/P3_XADDER/Xa13/Xyb2/M12_g N_VDD_XADDER/Xa13/Xyb2/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa0/M1 N_XCSA/XDFFA0/P001_XCSA/Xdffa0/M1_d
+ N_XCSA/LV3_C[1]_XCSA/Xdffa0/M1_g N_VDD_XCSA/Xdffa0/M1_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel20/M10 N_XBOOTH/XSEL20/B_XBOOTH/Xsel20/M10_d
+ N_XBOOTH/XSEL20/N002_XBOOTH/Xsel20/M10_g N_VDD_XBOOTH/Xsel20/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel10/M10 N_XBOOTH/XSEL10/B_XBOOTH/Xsel10/M10_d
+ N_XBOOTH/XSEL10/N002_XBOOTH/Xsel10/M10_g N_VDD_XBOOTH/Xsel10/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel00/M10 N_XBOOTH/XSEL00/B_XBOOTH/Xsel00/M10_d
+ N_XBOOTH/XSEL00/N002_XBOOTH/Xsel00/M10_g N_VDD_XBOOTH/Xsel00/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa13/M1 N_XCSA/XDFFA13/P001_XCSA/Xdffa13/M1_d
+ N_XCSA/LV3_S[1]_XCSA/Xdffa13/M1_g N_VDD_XCSA/Xdffa13/M1_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXADDER/Xa23/Xao2/M35 N_XADDER/XA23/XAO2/N007_XADDER/Xa23/Xao2/M35_d
+ N_XADDER/GG3_XADDER/Xa23/Xao2/M35_g N_VDD_XADDER/Xa23/Xao2/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXCSA/X_LV2_HA1/M10 N_XCSA/X_LV2_HA1/N001_XCSA/X_LV2_HA1/M10_d
+ N_A_D[3]_XCSA/X_LV2_HA1/M10_g N_VDD_XCSA/X_LV2_HA1/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA1/X_xor/M5 N_XCSA/X_LV2_HA1/X_XOR/N001_XCSA/X_LV2_HA1/X_xor/M5_d
+ N_A_D[3]_XCSA/X_LV2_HA1/X_xor/M5_g N_VDD_XCSA/X_LV2_HA1/X_xor/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXADDER/Xa04/Xrb2/M4 N_XADDER/P3_XADDER/Xa04/Xrb2/M4_d
+ N_XADDER/XA04/XRB2/N002_XADDER/Xa04/Xrb2/M4_g N_VDD_XADDER/Xa04/Xrb2/M4_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa0/M2 N_XCSA/XDFFA0/N0_XCSA/Xdffa0/M2_d N_CLK_XCSA/Xdffa0/M2_g
+ N_XCSA/XDFFA0/P001_XCSA/Xdffa0/M2_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa13/M2 N_XCSA/XDFFA13/N0_XCSA/Xdffa13/M2_d N_CLK_XCSA/Xdffa13/M2_g
+ N_XCSA/XDFFA13/P001_XCSA/Xdffa13/M2_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa13/Xyb2/M11 N_XADDER/XA13/XYB2/N003_XADDER/Xa13/Xyb2/M11_d
+ N_XADDER/G2_XADDER/Xa13/Xyb2/M11_g N_VDD_XADDER/Xa13/Xyb2/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mXCSA/X_LV2_HA1/X_xor/M6 N_XCSA/X_LV2_HA1/X_XOR/N002_XCSA/X_LV2_HA1/X_xor/M6_d
+ N_XCSA/LV1_S[2]_XCSA/X_LV2_HA1/X_xor/M6_g
+ N_XCSA/X_LV2_HA1/X_XOR/N001_XCSA/X_LV2_HA1/X_xor/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV3_HA0/X_xor/M6 N_XCSA/X_LV3_HA0/X_XOR/N001_XCSA/X_LV3_HA0/X_xor/M6_d
+ N_XCSA/LV2_S[0]_XCSA/X_LV3_HA0/X_xor/M6_g N_VDD_XCSA/X_LV3_HA0/X_xor/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV3_HA0/M9 N_XCSA/X_LV3_HA0/N001_XCSA/X_LV3_HA0/M9_d
+ N_XCSA/LV2_S[0]_XCSA/X_LV3_HA0/M9_g N_VDD_XCSA/X_LV3_HA0/M9_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXADDER/Xa23/Xao2/Xor1/M15 N_VDD_XADDER/Xa23/Xao2/Xor1/M15_d
+ N_XADDER/XA23/XAO2/N008_XADDER/Xa23/Xao2/Xor1/M15_g
+ N_XADDER/GGG3_XADDER/Xa23/Xao2/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mXCSA/X_LV2_HA1/M9 N_XCSA/X_LV2_HA1/N001_XCSA/X_LV2_HA1/M9_d
+ N_XCSA/LV1_S[2]_XCSA/X_LV2_HA1/M9_g N_VDD_XCSA/X_LV2_HA1/M9_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xdffb0/M4 N_XBOOTH/XDFFB0/N1_XBOOTH/Xdffb0/M4_d N_CLK_XBOOTH/Xdffb0/M4_g
+ N_VDD_XBOOTH/Xdffb0/M4_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07
+ AD=2.695e-13 AS=1.485e-13 PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_HA0/X_xor/M5 N_XCSA/X_LV3_HA0/X_XOR/N002_XCSA/X_LV3_HA0/X_xor/M5_d
+ N_CACC[0]_XCSA/X_LV3_HA0/X_xor/M5_g
+ N_XCSA/X_LV3_HA0/X_XOR/N001_XCSA/X_LV3_HA0/X_xor/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV1_HA0/M10 N_XCSA/X_LV1_HA0/N001_XCSA/X_LV1_HA0/M10_d
+ N_PP1[0]_XCSA/X_LV1_HA0/M10_g N_VDD_XCSA/X_LV1_HA0/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mX02/xd24/M4 N_X02/XD24/N1_X02/xd24/M4_d N_CLK_X02/xd24/M4_g N_VDD_X02/xd24/M4_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_HA0/M10 N_XCSA/X_LV3_HA0/N001_XCSA/X_LV3_HA0/M10_d
+ N_CACC[0]_XCSA/X_LV3_HA0/M10_g N_VDD_XCSA/X_LV3_HA0/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_HA0/X_xor/M5 N_XCSA/X_LV1_HA0/X_XOR/N002_XCSA/X_LV1_HA0/X_xor/M5_d
+ N_PP1[0]_XCSA/X_LV1_HA0/X_xor/M5_g
+ N_XCSA/X_LV1_HA0/X_XOR/N001_XCSA/X_LV1_HA0/X_xor/M5_s N_VDD_XBOOTH/Xdffa4/M1_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel20/M16 N_XBOOTH/XSEL20/N003_XBOOTH/Xsel20/M16_d
+ N_A_D[5]_XBOOTH/Xsel20/M16_g N_VDD_XBOOTH/Xsel20/M16_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel10/M16 N_XBOOTH/XSEL10/N003_XBOOTH/Xsel10/M16_d
+ N_A_D[3]_XBOOTH/Xsel10/M16_g N_VDD_XBOOTH/Xsel10/M16_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel00/M16 N_XBOOTH/XSEL00/N003_XBOOTH/Xsel00/M16_d
+ N_A_D[1]_XBOOTH/Xsel00/M16_g N_VDD_XBOOTH/Xsel00/M16_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xdffb0/M7 N_XBOOTH/XDFFB0/N3_XBOOTH/Xdffb0/M7_d
+ N_XBOOTH/XDFFB0/N1_XBOOTH/Xdffb0/M7_g N_VDD_XBOOTH/Xdffb0/M7_s
+ N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXADDER/Xa04/Xrb2/M5 N_XADDER/XA04/XRB2/N001_XADDER/Xa04/Xrb2/M5_d
+ N_C[3]_XADDER/Xa04/Xrb2/M5_g N_VDD_XADDER/Xa04/Xrb2/M5_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.904e-13
+ PD=2.8e-07 PS=1.76e-06
mXCSA/X_LV1_HA0/X_xor/M6 N_XCSA/X_LV1_HA0/X_XOR/N001_XCSA/X_LV1_HA0/X_xor/M6_d
+ N_PP0[2]_XCSA/X_LV1_HA0/X_xor/M6_g N_VDD_XCSA/X_LV1_HA0/X_xor/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV1_HA0/M9 N_XCSA/X_LV1_HA0/N001_XCSA/X_LV1_HA0/M9_d
+ N_PP0[2]_XCSA/X_LV1_HA0/M9_g N_VDD_XCSA/X_LV1_HA0/M9_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/Xdffa0/M4 N_XCSA/XDFFA0/N1_XCSA/Xdffa0/M4_d N_CLK_XCSA/Xdffa0/M4_g
+ N_VDD_XCSA/Xdffa0/M4_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa13/M4 N_XCSA/XDFFA13/N1_XCSA/Xdffa13/M4_d N_CLK_XCSA/Xdffa13/M4_g
+ N_VDD_XCSA/Xdffa13/M4_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mX02/xd24/M7 N_X02/XD24/N3_X02/xd24/M7_d N_X02/XD24/N1_X02/xd24/M7_g
+ N_VDD_X02/xd24/M7_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXADDER/Xa13/Xyb2/Xand1/M15 N_VDD_XADDER/Xa13/Xyb2/Xand1/M15_d
+ N_XADDER/XA13/XYB2/N003_XADDER/Xa13/Xyb2/Xand1/M15_g
+ N_XADDER/XA13/T1_XADDER/Xa13/Xyb2/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel20/M15 N_XBOOTH/XSEL20/N004_XBOOTH/Xsel20/M15_d
+ N_XBOOTH/XSEL20/B_XBOOTH/Xsel20/M15_g N_XBOOTH/XSEL20/N003_XBOOTH/Xsel20/M15_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel10/M15 N_XBOOTH/XSEL10/N004_XBOOTH/Xsel10/M15_d
+ N_XBOOTH/XSEL10/B_XBOOTH/Xsel10/M15_g N_XBOOTH/XSEL10/N003_XBOOTH/Xsel10/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel00/M15 N_XBOOTH/XSEL00/N004_XBOOTH/Xsel00/M15_d
+ N_XBOOTH/XSEL00/B_XBOOTH/Xsel00/M15_g N_XBOOTH/XSEL00/N003_XBOOTH/Xsel00/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV2_HA1/M13 N_XCSA/LV2_C[3]_XCSA/X_LV2_HA1/M13_d
+ N_XCSA/X_LV2_HA1/N001_XCSA/X_LV2_HA1/M13_g N_VDD_XCSA/X_LV2_HA1/M13_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA1/X_xor/M4 N_XCSA/LV2_S[2]_XCSA/X_LV2_HA1/X_xor/M4_d
+ N_XCSA/X_LV2_HA1/X_XOR/N002_XCSA/X_LV2_HA1/X_xor/M4_g
+ N_VDD_XCSA/X_LV2_HA1/X_xor/M4_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa04/Xrb2/M6 N_XADDER/XA04/XRB2/N002_XADDER/Xa04/Xrb2/M6_d
+ N_S[3]_XADDER/Xa04/Xrb2/M6_g N_XADDER/XA04/XRB2/N001_XADDER/Xa04/Xrb2/M6_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa0/M7 N_XCSA/XDFFA0/N3_XCSA/Xdffa0/M7_d
+ N_XCSA/XDFFA0/N1_XCSA/Xdffa0/M7_g N_VDD_XCSA/Xdffa0/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa13/M7 N_XCSA/XDFFA13/N3_XCSA/Xdffa13/M7_d
+ N_XCSA/XDFFA13/N1_XCSA/Xdffa13/M7_g N_VDD_XCSA/Xdffa13/M7_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa55/Xao1/M11 N_XADDER/XA55/XAO1/N003_XADDER/Xa55/Xao1/M11_d
+ N_XADDER/GGG3_XADDER/Xa55/Xao1/M11_g N_VDD_XADDER/Xa55/Xao1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.474e-13
+ PD=1.42e-06 PS=6.7e-07
mXCSA/X_LV3_HA0/X_xor/M4 N_XCSA/LV3_S[0]_XCSA/X_LV3_HA0/X_xor/M4_d
+ N_XCSA/X_LV3_HA0/X_XOR/N002_XCSA/X_LV3_HA0/X_xor/M4_g
+ N_VDD_XCSA/X_LV3_HA0/X_xor/M4_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_HA0/M13 N_XCSA/LV3_C[1]_XCSA/X_LV3_HA0/M13_d
+ N_XCSA/X_LV3_HA0/N001_XCSA/X_LV3_HA0/M13_g N_VDD_XCSA/X_LV3_HA0/M13_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xdffb0/M10 N_XBOOTH/B_D[0]_XBOOTH/Xdffb0/M10_d
+ N_XBOOTH/XDFFB0/N3_XBOOTH/Xdffb0/M10_g N_VDD_XBOOTH/Xdffb0/M10_s
+ N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mX02/xd24/M10 N_OUT[3]_X02/xd24/M10_d N_X02/XD24/N3_X02/xd24/M10_g
+ N_VDD_X02/xd24/M10_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel20/M14 N_PP2[0]_XBOOTH/Xsel20/M14_d
+ N_XBOOTH/XSEL20/N004_XBOOTH/Xsel20/M14_g N_VDD_XBOOTH/Xsel20/M14_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel10/M14 N_PP1[0]_XBOOTH/Xsel10/M14_d
+ N_XBOOTH/XSEL10/N004_XBOOTH/Xsel10/M14_g N_VDD_XBOOTH/Xsel10/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel00/M14 N_PP0[0]_XBOOTH/Xsel00/M14_d
+ N_XBOOTH/XSEL00/N004_XBOOTH/Xsel00/M14_g N_VDD_XBOOTH/Xsel00/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa55/Xao1/M12 N_XADDER/XA55/XAO1/N003_XADDER/Xa55/Xao1/M12_d
+ N_XADDER/PP5_XADDER/Xa55/Xao1/M12_g N_VDD_XADDER/Xa55/Xao1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.288e-13 AS=1.474e-13
+ PD=1.48e-06 PS=6.7e-07
mXADDER/Xa13/Xyb3/M36 N_XADDER/XA13/XYB3/N008_XADDER/Xa13/Xyb3/M36_d
+ N_XADDER/XA13/T1_XADDER/Xa13/Xyb3/M36_g
+ N_XADDER/XA13/XYB3/N007_XADDER/Xa13/Xyb3/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXADDER/Xa04/Xrb1/M12 N_XADDER/XA04/XRB1/N003_XADDER/Xa04/Xrb1/M12_d
+ N_S[3]_XADDER/Xa04/Xrb1/M12_g N_VDD_XADDER/Xa04/Xrb1/M12_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa0/M10 N_C[1]_XCSA/Xdffa0/M10_d N_XCSA/XDFFA0/N3_XCSA/Xdffa0/M10_g
+ N_VDD_XCSA/Xdffa0/M10_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa13/M10 N_S[1]_XCSA/Xdffa13/M10_d N_XCSA/XDFFA13/N3_XCSA/Xdffa13/M10_g
+ N_VDD_XCSA/Xdffa13/M10_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_HA1/X_xor/M4 N_XCSA/LV1_S[3]_XCSA/X_LV1_HA1/X_xor/M4_d
+ N_XCSA/X_LV1_HA1/X_XOR/N002_XCSA/X_LV1_HA1/X_xor/M4_g
+ N_VDD_XCSA/X_LV1_HA1/X_xor/M4_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_HA1/M13 N_XCSA/LV1_C[4]_XCSA/X_LV1_HA1/M13_d
+ N_XCSA/X_LV1_HA1/N001_XCSA/X_LV1_HA1/M13_g N_VDD_XCSA/X_LV1_HA1/M13_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa13/Xyb3/M35 N_XADDER/XA13/XYB3/N007_XADDER/Xa13/Xyb3/M35_d
+ N_XADDER/G3_XADDER/Xa13/Xyb3/M35_g N_VDD_XADDER/Xa13/Xyb3/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXCSA/X_LV2_HA2/M9 N_XCSA/X_LV2_HA2/N001_XCSA/X_LV2_HA2/M9_d
+ N_XCSA/LV1_C[3]_XCSA/X_LV2_HA2/M9_g N_VDD_XCSA/X_LV2_HA2/M9_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA2/X_xor/M6 N_XCSA/X_LV2_HA2/X_XOR/N001_XCSA/X_LV2_HA2/X_xor/M6_d
+ N_XCSA/LV1_C[3]_XCSA/X_LV2_HA2/X_xor/M6_g N_VDD_XCSA/X_LV2_HA2/X_xor/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXADDER/Xa04/Xrb1/M11 N_XADDER/XA04/XRB1/N003_XADDER/Xa04/Xrb1/M11_d
+ N_C[3]_XADDER/Xa04/Xrb1/M11_g N_VDD_XADDER/Xa04/Xrb1/M11_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA0/M27 N_XCSA/LV3_S[1]_XCSA/X_LV3_FA0/M27_d
+ N_XCSA/X_LV3_FA0/_SUM_XCSA/X_LV3_FA0/M27_g N_VDD_XCSA/X_LV3_FA0/M27_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mX02/xd25/M1 N_X02/XD25/P001_X02/xd25/M1_d N_OUT1[4]_X02/xd25/M1_g
+ N_VDD_X02/xd25/M1_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14
+ AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXADDER/Xa55/Xao1/Xand1/M15 N_VDD_XADDER/Xa55/Xao1/Xand1/M15_d
+ N_XADDER/XA55/XAO1/N003_XADDER/Xa55/Xao1/Xand1/M15_g
+ N_XADDER/XA55/OUT1_XADDER/Xa55/Xao1/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA2/X_xor/M5 N_XCSA/X_LV2_HA2/X_XOR/N002_XCSA/X_LV2_HA2/X_xor/M5_d
+ N_XCSA/LV1_S[3]_XCSA/X_LV2_HA2/X_xor/M5_g
+ N_XCSA/X_LV2_HA2/X_XOR/N001_XCSA/X_LV2_HA2/X_xor/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa13/Xyb3/Xor1/M15 N_VDD_XADDER/Xa13/Xyb3/Xor1/M15_d
+ N_XADDER/XA13/XYB3/N008_XADDER/Xa13/Xyb3/Xor1/M15_g
+ N_XADDER/GG3_XADDER/Xa13/Xyb3/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mXCSA/X_LV2_HA2/M10 N_XCSA/X_LV2_HA2/N001_XCSA/X_LV2_HA2/M10_d
+ N_XCSA/LV1_S[3]_XCSA/X_LV2_HA2/M10_g N_VDD_XCSA/X_LV2_HA2/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mX02/xd25/M2 N_X02/XD25/N0_X02/xd25/M2_d N_CLK_X02/xd25/M2_g
+ N_X02/XD25/P001_X02/xd25/M2_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa1/M1 N_XCSA/XDFFA1/P001_XCSA/Xdffa1/M1_d
+ N_XCSA/LV3_C[2]_XCSA/Xdffa1/M1_g N_VDD_XCSA/Xdffa1/M1_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa14/M1 N_XCSA/XDFFA14/P001_XCSA/Xdffa14/M1_d
+ N_XCSA/LV3_S[2]_XCSA/Xdffa14/M1_g N_VDD_XCSA/Xdffa14/M1_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV3_FA0/M28 N_XCSA/LV3_C[2]_XCSA/X_LV3_FA0/M28_d
+ N_XCSA/X_LV3_FA0/_COUT_XCSA/X_LV3_FA0/M28_g N_VDD_XCSA/X_LV3_FA0/M28_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXCSA/X_LV1_HA1/M10 N_XCSA/X_LV1_HA1/N001_XCSA/X_LV1_HA1/M10_d
+ N_PP1[1]_XCSA/X_LV1_HA1/M10_g N_VDD_XCSA/X_LV1_HA1/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel21/M8 N_XBOOTH/XSEL21/N002_XBOOTH/Xsel21/M8_d
+ N_XBOOTH/B_D[0]_XBOOTH/Xsel21/M8_g N_noxref_1548_XBOOTH/Xsel21/M8_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel11/M8 N_XBOOTH/XSEL11/N002_XBOOTH/Xsel11/M8_d
+ N_XBOOTH/B_D[0]_XBOOTH/Xsel11/M8_g N_noxref_1549_XBOOTH/Xsel11/M8_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel01/M8 N_XBOOTH/XSEL01/N002_XBOOTH/Xsel01/M8_d
+ N_XBOOTH/B_D[0]_XBOOTH/Xsel01/M8_g N_noxref_1550_XBOOTH/Xsel01/M8_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_HA1/X_xor/M5 N_XCSA/X_LV1_HA1/X_XOR/N002_XCSA/X_LV1_HA1/X_xor/M5_d
+ N_PP1[1]_XCSA/X_LV1_HA1/X_xor/M5_g
+ N_XCSA/X_LV1_HA1/X_XOR/N001_XCSA/X_LV1_HA1/X_xor/M5_s N_VDD_XBOOTH/Xdffa4/M1_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa1/M2 N_XCSA/XDFFA1/N0_XCSA/Xdffa1/M2_d N_CLK_XCSA/Xdffa1/M2_g
+ N_XCSA/XDFFA1/P001_XCSA/Xdffa1/M2_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa14/M2 N_XCSA/XDFFA14/N0_XCSA/Xdffa14/M2_d N_CLK_XCSA/Xdffa14/M2_g
+ N_XCSA/XDFFA14/P001_XCSA/Xdffa14/M2_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa04/Xrb1/Xand1/M15 N_VDD_XADDER/Xa04/Xrb1/Xand1/M15_d
+ N_XADDER/XA04/XRB1/N003_XADDER/Xa04/Xrb1/Xand1/M15_g
+ N_XADDER/G3_XADDER/Xa04/Xrb1/Xand1/M15_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA0/M9 N_XCSA/X_LV3_FA0/_SUM_XCSA/X_LV3_FA0/M9_d
+ N_XCSA/X_LV3_FA0/_COUT_XCSA/X_LV3_FA0/M9_g
+ N_XCSA/X_LV3_FA0/N002_XCSA/X_LV3_FA0/M9_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXCSA/X_LV1_HA1/X_xor/M6 N_XCSA/X_LV1_HA1/X_XOR/N001_XCSA/X_LV1_HA1/X_xor/M6_d
+ N_PP0[3]_XCSA/X_LV1_HA1/X_xor/M6_g N_VDD_XCSA/X_LV1_HA1/X_xor/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV1_HA1/M9 N_XCSA/X_LV1_HA1/N001_XCSA/X_LV1_HA1/M9_d
+ N_PP0[3]_XCSA/X_LV1_HA1/M9_g N_VDD_XCSA/X_LV1_HA1/M9_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXBOOTH/Xsel21/M6 N_XBOOTH/XSEL21/N002_XBOOTH/Xsel21/M6_d
+ N_XBOOTH/D2_XBOOTH/Xsel21/M6_g N_noxref_1548_XBOOTH/Xsel21/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel11/M6 N_XBOOTH/XSEL11/N002_XBOOTH/Xsel11/M6_d
+ N_XBOOTH/D1_XBOOTH/Xsel11/M6_g N_noxref_1549_XBOOTH/Xsel11/M6_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel01/M6 N_XBOOTH/XSEL01/N002_XBOOTH/Xsel01/M6_d
+ N_XBOOTH/D0_XBOOTH/Xsel01/M6_g N_noxref_1550_XBOOTH/Xsel01/M6_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXADDER/Xa55/Xao2/M36 N_XADDER/XA55/XAO2/N008_XADDER/Xa55/Xao2/M36_d
+ N_XADDER/XA55/OUT1_XADDER/Xa55/Xao2/M36_g
+ N_XADDER/XA55/XAO2/N007_XADDER/Xa55/Xao2/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXCSA/X_LV2_HA2/M13 N_XCSA/LV2_C[4]_XCSA/X_LV2_HA2/M13_d
+ N_XCSA/X_LV2_HA2/N001_XCSA/X_LV2_HA2/M13_g N_VDD_XCSA/X_LV2_HA2/M13_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA2/X_xor/M4 N_XCSA/LV2_S[3]_XCSA/X_LV2_HA2/X_xor/M4_d
+ N_XCSA/X_LV2_HA2/X_XOR/N002_XCSA/X_LV2_HA2/X_xor/M4_g
+ N_VDD_XCSA/X_LV2_HA2/X_xor/M4_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd25/M4 N_X02/XD25/N1_X02/xd25/M4_d N_CLK_X02/xd25/M4_g N_VDD_X02/xd25/M4_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa15/Xyb1/Xand1/M15 N_VDD_XADDER/Xa15/Xyb1/Xand1/M15_d
+ N_XADDER/XA15/XYB1/N003_XADDER/Xa15/Xyb1/Xand1/M15_g
+ N_XADDER/PP5_XADDER/Xa15/Xyb1/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA0/M5 N_XCSA/X_LV3_FA0/_COUT_XCSA/X_LV3_FA0/M5_d
+ N_CACC[1]_XCSA/X_LV3_FA0/M5_g N_XCSA/X_LV3_FA0/N001_XCSA/X_LV3_FA0/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA0/M12 N_XCSA/X_LV3_FA0/_SUM_XCSA/X_LV3_FA0/M12_d
+ N_CACC[1]_XCSA/X_LV3_FA0/M12_g N_XCSA/X_LV3_FA0/P003_XCSA/X_LV3_FA0/M12_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA0/M6 N_XCSA/X_LV3_FA0/N002_XCSA/X_LV3_FA0/M6_d
+ N_CACC[1]_XCSA/X_LV3_FA0/M6_g N_VDD_XCSA/X_LV3_FA0/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXBOOTH/Xsel21/M7 N_noxref_1548_XBOOTH/Xsel21/M7_d
+ N_XBOOTH/S2_XBOOTH/Xsel21/M7_g N_VDD_XBOOTH/Xsel21/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel11/M7 N_noxref_1549_XBOOTH/Xsel11/M7_d
+ N_XBOOTH/S1_XBOOTH/Xsel11/M7_g N_VDD_XBOOTH/Xsel11/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel01/M7 N_noxref_1550_XBOOTH/Xsel01/M7_d
+ N_XBOOTH/S0_XBOOTH/Xsel01/M7_g N_VDD_XBOOTH/Xsel01/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXADDER/Xa55/Xao2/M35 N_XADDER/XA55/XAO2/N007_XADDER/Xa55/Xao2/M35_d
+ N_XADDER/GG5_XADDER/Xa55/Xao2/M35_g N_VDD_XADDER/Xa55/Xao2/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXCSA/Xdffa1/M4 N_XCSA/XDFFA1/N1_XCSA/Xdffa1/M4_d N_CLK_XCSA/Xdffa1/M4_g
+ N_VDD_XCSA/Xdffa1/M4_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa14/M4 N_XCSA/XDFFA14/N1_XCSA/Xdffa14/M4_d N_CLK_XCSA/Xdffa14/M4_g
+ N_VDD_XCSA/Xdffa14/M4_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mX02/xd25/M7 N_X02/XD25/N3_X02/xd25/M7_d N_X02/XD25/N1_X02/xd25/M7_g
+ N_VDD_X02/xd25/M7_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXADDER/Xa05/Xrb2/M4 N_XADDER/P4_XADDER/Xa05/Xrb2/M4_d
+ N_XADDER/XA05/XRB2/N002_XADDER/Xa05/Xrb2/M4_g N_VDD_XADDER/Xa05/Xrb2/M4_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xdffb1/M1 N_XBOOTH/XDFFB1/P001_XBOOTH/Xdffb1/M1_d
+ N_B[1]_XBOOTH/Xdffb1/M1_g N_VDD_XBOOTH/Xdffb1/M1_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=7.7e-14 AS=2.695e-13 PD=2.8e-07 PS=1.53e-06
mXCSA/X_LV3_FA0/M4 N_XCSA/X_LV3_FA0/N001_XCSA/X_LV3_FA0/M4_d
+ N_PP0[1]_XCSA/X_LV3_FA0/M4_g N_VDD_XCSA/X_LV3_FA0/M4_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA0/M2 N_XCSA/X_LV3_FA0/_COUT_XCSA/X_LV3_FA0/M2_d
+ N_PP0[1]_XCSA/X_LV3_FA0/M2_g N_XCSA/X_LV3_FA0/P001_XCSA/X_LV3_FA0/M2_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA0/M11 N_XCSA/X_LV3_FA0/P003_XCSA/X_LV3_FA0/M11_d
+ N_PP0[1]_XCSA/X_LV3_FA0/M11_g N_XCSA/X_LV3_FA0/P002_XCSA/X_LV3_FA0/M11_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA0/M8 N_XCSA/X_LV3_FA0/N002_XCSA/X_LV3_FA0/M8_d
+ N_PP0[1]_XCSA/X_LV3_FA0/M8_g N_VDD_XCSA/X_LV3_FA0/M8_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mXBOOTH/Xsel21/M9 N_noxref_1548_XBOOTH/Xsel21/M9_d
+ N_XBOOTH/B_D[1]_XBOOTH/Xsel21/M9_g N_VDD_XBOOTH/Xsel21/M9_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel11/M9 N_noxref_1549_XBOOTH/Xsel11/M9_d
+ N_XBOOTH/B_D[1]_XBOOTH/Xsel11/M9_g N_VDD_XBOOTH/Xsel11/M9_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel01/M9 N_noxref_1550_XBOOTH/Xsel01/M9_d
+ N_XBOOTH/B_D[1]_XBOOTH/Xsel01/M9_g N_VDD_XBOOTH/Xsel01/M9_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa55/Xao2/Xor1/M15 N_VDD_XADDER/Xa55/Xao2/Xor1/M15_d
+ N_XADDER/XA55/XAO2/N008_XADDER/Xa55/Xao2/Xor1/M15_g
+ N_XADDER/GX5[0]_XADDER/Xa55/Xao2/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mXBOOTH/Xdffb1/M2 N_XBOOTH/XDFFB1/N0_XBOOTH/Xdffb1/M2_d N_CLK_XBOOTH/Xdffb1/M2_g
+ N_XBOOTH/XDFFB1/P001_XBOOTH/Xdffb1/M2_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=7.7e-14 PD=1.53e-06 PS=2.8e-07
mXCSA/Xdffa1/M7 N_XCSA/XDFFA1/N3_XCSA/Xdffa1/M7_d
+ N_XCSA/XDFFA1/N1_XCSA/Xdffa1/M7_g N_VDD_XCSA/Xdffa1/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa14/M7 N_XCSA/XDFFA14/N3_XCSA/Xdffa14/M7_d
+ N_XCSA/XDFFA14/N1_XCSA/Xdffa14/M7_g N_VDD_XCSA/Xdffa14/M7_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA0/M3 N_XCSA/X_LV3_FA0/N001_XCSA/X_LV3_FA0/M3_d
+ N_XCSA/LV2_C[1]_XCSA/X_LV3_FA0/M3_g N_VDD_XCSA/X_LV3_FA0/M3_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA0/M1 N_XCSA/X_LV3_FA0/P001_XCSA/X_LV3_FA0/M1_d
+ N_XCSA/LV2_C[1]_XCSA/X_LV3_FA0/M1_g N_VDD_XCSA/X_LV3_FA0/M1_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA0/M10 N_XCSA/X_LV3_FA0/P002_XCSA/X_LV3_FA0/M10_d
+ N_XCSA/LV2_C[1]_XCSA/X_LV3_FA0/M10_g N_VDD_XCSA/X_LV3_FA0/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA0/M7 N_XCSA/X_LV3_FA0/N002_XCSA/X_LV3_FA0/M7_d
+ N_XCSA/LV2_C[1]_XCSA/X_LV3_FA0/M7_g N_VDD_XCSA/X_LV3_FA0/M7_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXADDER/Xa15/Xyb1/M11 N_XADDER/XA15/XYB1/N003_XADDER/Xa15/Xyb1/M11_d
+ N_XADDER/P4_XADDER/Xa15/Xyb1/M11_g N_VDD_XADDER/Xa15/Xyb1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mXBOOTH/Xsel21/M10 N_XBOOTH/XSEL21/B_XBOOTH/Xsel21/M10_d
+ N_XBOOTH/XSEL21/N002_XBOOTH/Xsel21/M10_g N_VDD_XBOOTH/Xsel21/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel11/M10 N_XBOOTH/XSEL11/B_XBOOTH/Xsel11/M10_d
+ N_XBOOTH/XSEL11/N002_XBOOTH/Xsel11/M10_g N_VDD_XBOOTH/Xsel11/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel01/M10 N_XBOOTH/XSEL01/B_XBOOTH/Xsel01/M10_d
+ N_XBOOTH/XSEL01/N002_XBOOTH/Xsel01/M10_g N_VDD_XBOOTH/Xsel01/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA0/M3 N_XCSA/X_LV1_FA0/N001_XCSA/X_LV1_FA0/M3_d
+ N_PP0[4]_XCSA/X_LV1_FA0/M3_g N_VDD_XCSA/X_LV1_FA0/M3_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV1_FA0/M1 N_XCSA/X_LV1_FA0/P001_XCSA/X_LV1_FA0/M1_d
+ N_PP0[4]_XCSA/X_LV1_FA0/M1_g N_VDD_XCSA/X_LV1_FA0/M1_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV1_FA0/M10 N_XCSA/X_LV1_FA0/P002_XCSA/X_LV1_FA0/M10_d
+ N_PP0[4]_XCSA/X_LV1_FA0/M10_g N_VDD_XCSA/X_LV1_FA0/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV1_FA0/M7 N_XCSA/X_LV1_FA0/N002_XCSA/X_LV1_FA0/M7_d
+ N_PP0[4]_XCSA/X_LV1_FA0/M7_g N_VDD_XCSA/X_LV1_FA0/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mX02/xd25/M10 N_OUT[4]_X02/xd25/M10_d N_X02/XD25/N3_X02/xd25/M10_g
+ N_VDD_X02/xd25/M10_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_FA0/M7 N_XCSA/X_LV2_FA0/N002_XCSA/X_LV2_FA0/M7_d
+ N_XCSA/LV1_C[4]_XCSA/X_LV2_FA0/M7_g N_VDD_XCSA/X_LV2_FA0/M7_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV2_FA0/M10 N_XCSA/X_LV2_FA0/P002_XCSA/X_LV2_FA0/M10_d
+ N_XCSA/LV1_C[4]_XCSA/X_LV2_FA0/M10_g N_VDD_XCSA/X_LV2_FA0/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV2_FA0/M1 N_XCSA/X_LV2_FA0/P001_XCSA/X_LV2_FA0/M1_d
+ N_XCSA/LV1_C[4]_XCSA/X_LV2_FA0/M1_g N_VDD_XCSA/X_LV2_FA0/M1_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV2_FA0/M3 N_XCSA/X_LV2_FA0/N001_XCSA/X_LV2_FA0/M3_d
+ N_XCSA/LV1_C[4]_XCSA/X_LV2_FA0/M3_g N_VDD_XCSA/X_LV2_FA0/M3_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXADDER/Xa05/Xrb2/M5 N_XADDER/XA05/XRB2/N001_XADDER/Xa05/Xrb2/M5_d
+ N_C[4]_XADDER/Xa05/Xrb2/M5_g N_VDD_XADDER/Xa05/Xrb2/M5_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.904e-13
+ PD=2.8e-07 PS=1.76e-06
mXADDER/Xa15/Xyb1/M12 N_XADDER/XA15/XYB1/N003_XADDER/Xa15/Xyb1/M12_d
+ N_XADDER/P5_XADDER/Xa15/Xyb1/M12_g N_VDD_XADDER/Xa15/Xyb1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xdffb1/M4 N_XBOOTH/XDFFB1/N1_XBOOTH/Xdffb1/M4_d N_CLK_XBOOTH/Xdffb1/M4_g
+ N_VDD_XBOOTH/Xdffb1/M4_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07
+ AD=2.695e-13 AS=1.485e-13 PD=1.53e-06 PS=5.4e-07
mXCSA/Xdffa1/M10 N_C[2]_XCSA/Xdffa1/M10_d N_XCSA/XDFFA1/N3_XCSA/Xdffa1/M10_g
+ N_VDD_XCSA/Xdffa1/M10_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa14/M10 N_S[2]_XCSA/Xdffa14/M10_d N_XCSA/XDFFA14/N3_XCSA/Xdffa14/M10_g
+ N_VDD_XCSA/Xdffa14/M10_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA0/M4 N_XCSA/X_LV1_FA0/N001_XCSA/X_LV1_FA0/M4_d
+ N_PP1[2]_XCSA/X_LV1_FA0/M4_g N_VDD_XCSA/X_LV1_FA0/M4_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA0/M2 N_XCSA/X_LV1_FA0/_COUT_XCSA/X_LV1_FA0/M2_d
+ N_PP1[2]_XCSA/X_LV1_FA0/M2_g N_XCSA/X_LV1_FA0/P001_XCSA/X_LV1_FA0/M2_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV1_FA0/M11 N_XCSA/X_LV1_FA0/P003_XCSA/X_LV1_FA0/M11_d
+ N_PP1[2]_XCSA/X_LV1_FA0/M11_g N_XCSA/X_LV1_FA0/P002_XCSA/X_LV1_FA0/M11_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA0/M8 N_XCSA/X_LV1_FA0/N002_XCSA/X_LV1_FA0/M8_d
+ N_PP1[2]_XCSA/X_LV1_FA0/M8_g N_VDD_XCSA/X_LV1_FA0/M8_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mXADDER/Xa05/Xrb2/M6 N_XADDER/XA05/XRB2/N002_XADDER/Xa05/Xrb2/M6_d
+ N_S[4]_XADDER/Xa05/Xrb2/M6_g N_XADDER/XA05/XRB2/N001_XADDER/Xa05/Xrb2/M6_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV2_FA0/M8 N_XCSA/X_LV2_FA0/N002_XCSA/X_LV2_FA0/M8_d
+ N_XCSA/LV1_S[4]_XCSA/X_LV2_FA0/M8_g N_VDD_XCSA/X_LV2_FA0/M8_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV2_FA0/M11 N_XCSA/X_LV2_FA0/P003_XCSA/X_LV2_FA0/M11_d
+ N_XCSA/LV1_S[4]_XCSA/X_LV2_FA0/M11_g
+ N_XCSA/X_LV2_FA0/P002_XCSA/X_LV2_FA0/M11_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV2_FA0/M2 N_XCSA/X_LV2_FA0/_COUT_XCSA/X_LV2_FA0/M2_d
+ N_XCSA/LV1_S[4]_XCSA/X_LV2_FA0/M2_g N_XCSA/X_LV2_FA0/P001_XCSA/X_LV2_FA0/M2_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV2_FA0/M4 N_XCSA/X_LV2_FA0/N001_XCSA/X_LV2_FA0/M4_d
+ N_XCSA/LV1_S[4]_XCSA/X_LV2_FA0/M4_g N_VDD_XCSA/X_LV2_FA0/M4_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXADDER/Xa64/Xao1/M11 N_XADDER/XA64/XAO1/N003_XADDER/Xa64/Xao1/M11_d
+ N_XADDER/GGG3_XADDER/Xa64/Xao1/M11_g N_VDD_XADDER/Xa64/Xao1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.474e-13
+ PD=1.42e-06 PS=6.7e-07
mXBOOTH/Xdffb1/M7 N_XBOOTH/XDFFB1/N3_XBOOTH/Xdffb1/M7_d
+ N_XBOOTH/XDFFB1/N1_XBOOTH/Xdffb1/M7_g N_VDD_XBOOTH/Xdffb1/M7_s
+ N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mX02/xd26/M1 N_X02/XD26/P001_X02/xd26/M1_d N_OUT1[5]_X02/xd26/M1_g
+ N_VDD_X02/xd26/M1_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14
+ AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV1_FA0/M5 N_XCSA/X_LV1_FA0/_COUT_XCSA/X_LV1_FA0/M5_d
+ N_PP2[0]_XCSA/X_LV1_FA0/M5_g N_XCSA/X_LV1_FA0/N001_XCSA/X_LV1_FA0/M5_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV1_FA0/M12 N_XCSA/X_LV1_FA0/_SUM_XCSA/X_LV1_FA0/M12_d
+ N_PP2[0]_XCSA/X_LV1_FA0/M12_g N_XCSA/X_LV1_FA0/P003_XCSA/X_LV1_FA0/M12_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV1_FA0/M6 N_XCSA/X_LV1_FA0/N002_XCSA/X_LV1_FA0/M6_d
+ N_PP2[0]_XCSA/X_LV1_FA0/M6_g N_VDD_XCSA/X_LV1_FA0/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV2_FA0/M6 N_XCSA/X_LV2_FA0/N002_XCSA/X_LV2_FA0/M6_d
+ N_A_D[5]_XCSA/X_LV2_FA0/M6_g N_VDD_XCSA/X_LV2_FA0/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV2_FA0/M12 N_XCSA/X_LV2_FA0/_SUM_XCSA/X_LV2_FA0/M12_d
+ N_A_D[5]_XCSA/X_LV2_FA0/M12_g N_XCSA/X_LV2_FA0/P003_XCSA/X_LV2_FA0/M12_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV2_FA0/M5 N_XCSA/X_LV2_FA0/_COUT_XCSA/X_LV2_FA0/M5_d
+ N_A_D[5]_XCSA/X_LV2_FA0/M5_g N_XCSA/X_LV2_FA0/N001_XCSA/X_LV2_FA0/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXBOOTH/Xsel21/M16 N_XBOOTH/XSEL21/N003_XBOOTH/Xsel21/M16_d
+ N_A_D[5]_XBOOTH/Xsel21/M16_g N_VDD_XBOOTH/Xsel21/M16_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel11/M16 N_XBOOTH/XSEL11/N003_XBOOTH/Xsel11/M16_d
+ N_A_D[3]_XBOOTH/Xsel11/M16_g N_VDD_XBOOTH/Xsel11/M16_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel01/M16 N_XBOOTH/XSEL01/N003_XBOOTH/Xsel01/M16_d
+ N_A_D[1]_XBOOTH/Xsel01/M16_g N_VDD_XBOOTH/Xsel01/M16_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV3_HA1/X_xor/M6 N_XCSA/X_LV3_HA1/X_XOR/N001_XCSA/X_LV3_HA1/X_xor/M6_d
+ N_XCSA/LV2_S[2]_XCSA/X_LV3_HA1/X_xor/M6_g N_VDD_XCSA/X_LV3_HA1/X_xor/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV3_HA1/M9 N_XCSA/X_LV3_HA1/N001_XCSA/X_LV3_HA1/M9_d
+ N_XCSA/LV2_S[2]_XCSA/X_LV3_HA1/M9_g N_VDD_XCSA/X_LV3_HA1/M9_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXADDER/Xa15/Xyb2/M12 N_XADDER/XA15/XYB2/N003_XADDER/Xa15/Xyb2/M12_d
+ N_XADDER/P5_XADDER/Xa15/Xyb2/M12_g N_VDD_XADDER/Xa15/Xyb2/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd26/M2 N_X02/XD26/N0_X02/xd26/M2_d N_CLK_X02/xd26/M2_g
+ N_X02/XD26/P001_X02/xd26/M2_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa64/Xao1/M12 N_XADDER/XA64/XAO1/N003_XADDER/Xa64/Xao1/M12_d
+ N_XADDER/P4_XADDER/Xa64/Xao1/M12_g N_VDD_XADDER/Xa64/Xao1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.288e-13 AS=1.474e-13
+ PD=1.48e-06 PS=6.7e-07
mXCSA/Xdffa2/M1 N_XCSA/XDFFA2/P001_XCSA/Xdffa2/M1_d
+ N_XCSA/LV3_C[3]_XCSA/Xdffa2/M1_g N_VDD_XCSA/Xdffa2/M1_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel21/M15 N_XBOOTH/XSEL21/N004_XBOOTH/Xsel21/M15_d
+ N_XBOOTH/XSEL21/B_XBOOTH/Xsel21/M15_g N_XBOOTH/XSEL21/N003_XBOOTH/Xsel21/M15_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel11/M15 N_XBOOTH/XSEL11/N004_XBOOTH/Xsel11/M15_d
+ N_XBOOTH/XSEL11/B_XBOOTH/Xsel11/M15_g N_XBOOTH/XSEL11/N003_XBOOTH/Xsel11/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel01/M15 N_XBOOTH/XSEL01/N004_XBOOTH/Xsel01/M15_d
+ N_XBOOTH/XSEL01/B_XBOOTH/Xsel01/M15_g N_XBOOTH/XSEL01/N003_XBOOTH/Xsel01/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa15/M1 N_XCSA/XDFFA15/P001_XCSA/Xdffa15/M1_d
+ N_XCSA/LV3_S[3]_XCSA/Xdffa15/M1_g N_VDD_XCSA/Xdffa15/M1_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV3_HA1/X_xor/M5 N_XCSA/X_LV3_HA1/X_XOR/N002_XCSA/X_LV3_HA1/X_xor/M5_d
+ N_CACC[2]_XCSA/X_LV3_HA1/X_xor/M5_g
+ N_XCSA/X_LV3_HA1/X_XOR/N001_XCSA/X_LV3_HA1/X_xor/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV1_FA0/M9 N_XCSA/X_LV1_FA0/_SUM_XCSA/X_LV1_FA0/M9_d
+ N_XCSA/X_LV1_FA0/_COUT_XCSA/X_LV1_FA0/M9_g
+ N_XCSA/X_LV1_FA0/N002_XCSA/X_LV1_FA0/M9_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXCSA/X_LV3_HA1/M10 N_XCSA/X_LV3_HA1/N001_XCSA/X_LV3_HA1/M10_d
+ N_CACC[2]_XCSA/X_LV3_HA1/M10_g N_VDD_XCSA/X_LV3_HA1/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa05/Xrb1/M12 N_XADDER/XA05/XRB1/N003_XADDER/Xa05/Xrb1/M12_d
+ N_S[4]_XADDER/Xa05/Xrb1/M12_g N_VDD_XADDER/Xa05/Xrb1/M12_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV2_FA0/M9 N_XCSA/X_LV2_FA0/_SUM_XCSA/X_LV2_FA0/M9_d
+ N_XCSA/X_LV2_FA0/_COUT_XCSA/X_LV2_FA0/M9_g
+ N_XCSA/X_LV2_FA0/N002_XCSA/X_LV2_FA0/M9_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXCSA/Xdffa2/M2 N_XCSA/XDFFA2/N0_XCSA/Xdffa2/M2_d N_CLK_XCSA/Xdffa2/M2_g
+ N_XCSA/XDFFA2/P001_XCSA/Xdffa2/M2_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa15/M2 N_XCSA/XDFFA15/N0_XCSA/Xdffa15/M2_d N_CLK_XCSA/Xdffa15/M2_g
+ N_XCSA/XDFFA15/P001_XCSA/Xdffa15/M2_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa15/Xyb2/M11 N_XADDER/XA15/XYB2/N003_XADDER/Xa15/Xyb2/M11_d
+ N_XADDER/G4_XADDER/Xa15/Xyb2/M11_g N_VDD_XADDER/Xa15/Xyb2/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mXBOOTH/Xdffb1/M10 N_XBOOTH/B_D[1]_XBOOTH/Xdffb1/M10_d
+ N_XBOOTH/XDFFB1/N3_XBOOTH/Xdffb1/M10_g N_VDD_XBOOTH/Xdffb1/M10_s
+ N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa75/M4 N_OUT1[5]_XADDER/Xa75/M4_d N_XADDER/XA75/N002_XADDER/Xa75/M4_g
+ N_VDD_XADDER/Xa75/M4_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA0/M28 N_XCSA/LV1_C[5]_XCSA/X_LV1_FA0/M28_d
+ N_XCSA/X_LV1_FA0/_COUT_XCSA/X_LV1_FA0/M28_g N_VDD_XCSA/X_LV1_FA0/M28_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXCSA/X_LV2_FA0/M28 N_XCSA/LV2_C[5]_XCSA/X_LV2_FA0/M28_d
+ N_XCSA/X_LV2_FA0/_COUT_XCSA/X_LV2_FA0/M28_g N_VDD_XCSA/X_LV2_FA0/M28_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa05/Xrb1/M11 N_XADDER/XA05/XRB1/N003_XADDER/Xa05/Xrb1/M11_d
+ N_C[4]_XADDER/Xa05/Xrb1/M11_g N_VDD_XADDER/Xa05/Xrb1/M11_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd26/M4 N_X02/XD26/N1_X02/xd26/M4_d N_CLK_X02/xd26/M4_g N_VDD_X02/xd26/M4_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel21/M14 N_PP2[1]_XBOOTH/Xsel21/M14_d
+ N_XBOOTH/XSEL21/N004_XBOOTH/Xsel21/M14_g N_VDD_XBOOTH/Xsel21/M14_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel11/M14 N_PP1[1]_XBOOTH/Xsel11/M14_d
+ N_XBOOTH/XSEL11/N004_XBOOTH/Xsel11/M14_g N_VDD_XBOOTH/Xsel11/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel01/M14 N_PP0[1]_XBOOTH/Xsel01/M14_d
+ N_XBOOTH/XSEL01/N004_XBOOTH/Xsel01/M14_g N_VDD_XBOOTH/Xsel01/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa64/Xao1/Xand1/M15 N_VDD_XADDER/Xa64/Xao1/Xand1/M15_d
+ N_XADDER/XA64/XAO1/N003_XADDER/Xa64/Xao1/Xand1/M15_g
+ N_XADDER/XA64/OUT1_XADDER/Xa64/Xao1/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA0/M27 N_XCSA/LV1_S[4]_XCSA/X_LV1_FA0/M27_d
+ N_XCSA/X_LV1_FA0/_SUM_XCSA/X_LV1_FA0/M27_g N_VDD_XCSA/X_LV1_FA0/M27_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXCSA/X_LV3_HA1/X_xor/M4 N_XCSA/LV3_S[2]_XCSA/X_LV3_HA1/X_xor/M4_d
+ N_XCSA/X_LV3_HA1/X_XOR/N002_XCSA/X_LV3_HA1/X_xor/M4_g
+ N_VDD_XCSA/X_LV3_HA1/X_xor/M4_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_HA1/M13 N_XCSA/LV3_C[3]_XCSA/X_LV3_HA1/M13_d
+ N_XCSA/X_LV3_HA1/N001_XCSA/X_LV3_HA1/M13_g N_VDD_XCSA/X_LV3_HA1/M13_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_FA0/M27 N_XCSA/LV2_S[4]_XCSA/X_LV2_FA0/M27_d
+ N_XCSA/X_LV2_FA0/_SUM_XCSA/X_LV2_FA0/M27_g N_VDD_XCSA/X_LV2_FA0/M27_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXCSA/Xdffa2/M4 N_XCSA/XDFFA2/N1_XCSA/Xdffa2/M4_d N_CLK_XCSA/Xdffa2/M4_g
+ N_VDD_XCSA/Xdffa2/M4_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa15/M4 N_XCSA/XDFFA15/N1_XCSA/Xdffa15/M4_d N_CLK_XCSA/Xdffa15/M4_g
+ N_VDD_XCSA/Xdffa15/M4_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mX02/xd26/M7 N_X02/XD26/N3_X02/xd26/M7_d N_X02/XD26/N1_X02/xd26/M7_g
+ N_VDD_X02/xd26/M7_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXADDER/Xa15/Xyb2/Xand1/M15 N_VDD_XADDER/Xa15/Xyb2/Xand1/M15_d
+ N_XADDER/XA15/XYB2/N003_XADDER/Xa15/Xyb2/Xand1/M15_g
+ N_XADDER/XA15/T1_XADDER/Xa15/Xyb2/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa05/Xrb1/Xand1/M15 N_VDD_XADDER/Xa05/Xrb1/Xand1/M15_d
+ N_XADDER/XA05/XRB1/N003_XADDER/Xa05/Xrb1/Xand1/M15_g
+ N_XADDER/G4_XADDER/Xa05/Xrb1/Xand1/M15_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa2/M7 N_XCSA/XDFFA2/N3_XCSA/Xdffa2/M7_d
+ N_XCSA/XDFFA2/N1_XCSA/Xdffa2/M7_g N_VDD_XCSA/Xdffa2/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa15/M7 N_XCSA/XDFFA15/N3_XCSA/Xdffa15/M7_d
+ N_XCSA/XDFFA15/N1_XCSA/Xdffa15/M7_g N_VDD_XCSA/Xdffa15/M7_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa75/M5 N_XADDER/XA75/N002_XADDER/Xa75/M5_d N_XADDER/P5_XADDER/Xa75/M5_g
+ N_XADDER/XA75/N001_XADDER/Xa75/M5_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=4.444e-13 AS=6.16e-14 PD=2.46e-06 PS=2.8e-07
mXADDER/Xa64/Xao2/M36 N_XADDER/XA64/XAO2/N008_XADDER/Xa64/Xao2/M36_d
+ N_XADDER/XA64/OUT1_XADDER/Xa64/Xao2/M36_g
+ N_XADDER/XA64/XAO2/N007_XADDER/Xa64/Xao2/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXADDER/Xa75/M6 N_XADDER/XA75/N001_XADDER/Xa75/M6_d
+ N_XADDER/GX6[1]_XADDER/Xa75/M6_g N_VDD_XADDER/Xa75/M6_s N_VDD_XADDER/Xa72/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mX02/xd26/M10 N_OUT[5]_X02/xd26/M10_d N_X02/XD26/N3_X02/xd26/M10_g
+ N_VDD_X02/xd26/M10_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel22/M8 N_XBOOTH/XSEL22/N002_XBOOTH/Xsel22/M8_d
+ N_XBOOTH/B_D[1]_XBOOTH/Xsel22/M8_g N_noxref_1594_XBOOTH/Xsel22/M8_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel12/M8 N_XBOOTH/XSEL12/N002_XBOOTH/Xsel12/M8_d
+ N_XBOOTH/B_D[1]_XBOOTH/Xsel12/M8_g N_noxref_1595_XBOOTH/Xsel12/M8_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel02/M8 N_XBOOTH/XSEL02/N002_XBOOTH/Xsel02/M8_d
+ N_XBOOTH/B_D[1]_XBOOTH/Xsel02/M8_g N_noxref_1596_XBOOTH/Xsel02/M8_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa64/Xao2/M35 N_XADDER/XA64/XAO2/N007_XADDER/Xa64/Xao2/M35_d
+ N_XADDER/G4_XADDER/Xa64/Xao2/M35_g N_VDD_XADDER/Xa64/Xao2/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXADDER/Xa15/Xyb3/M36 N_XADDER/XA15/XYB3/N008_XADDER/Xa15/Xyb3/M36_d
+ N_XADDER/XA15/T1_XADDER/Xa15/Xyb3/M36_g
+ N_XADDER/XA15/XYB3/N007_XADDER/Xa15/Xyb3/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXCSA/X_LV2_HA3/M9 N_XCSA/X_LV2_HA3/N001_XCSA/X_LV2_HA3/M9_d
+ N_XCSA/LV1_C[5]_XCSA/X_LV2_HA3/M9_g N_VDD_XCSA/X_LV2_HA3/M9_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA3/X_xor/M6 N_XCSA/X_LV2_HA3/X_XOR/N001_XCSA/X_LV2_HA3/X_xor/M6_d
+ N_XCSA/LV1_C[5]_XCSA/X_LV2_HA3/X_xor/M6_g N_VDD_XCSA/X_LV2_HA3/X_xor/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV3_FA1/M27 N_XCSA/LV3_S[3]_XCSA/X_LV3_FA1/M27_d
+ N_XCSA/X_LV3_FA1/_SUM_XCSA/X_LV3_FA1/M27_g N_VDD_XCSA/X_LV3_FA1/M27_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXCSA/X_LV1_FA1/M3 N_XCSA/X_LV1_FA1/N001_XCSA/X_LV1_FA1/M3_d
+ N_PP0[5]_XCSA/X_LV1_FA1/M3_g N_VDD_XCSA/X_LV1_FA1/M3_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV1_FA1/M1 N_XCSA/X_LV1_FA1/P001_XCSA/X_LV1_FA1/M1_d
+ N_PP0[5]_XCSA/X_LV1_FA1/M1_g N_VDD_XCSA/X_LV1_FA1/M1_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV1_FA1/M10 N_XCSA/X_LV1_FA1/P002_XCSA/X_LV1_FA1/M10_d
+ N_PP0[5]_XCSA/X_LV1_FA1/M10_g N_VDD_XCSA/X_LV1_FA1/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV1_FA1/M7 N_XCSA/X_LV1_FA1/N002_XCSA/X_LV1_FA1/M7_d
+ N_PP0[5]_XCSA/X_LV1_FA1/M7_g N_VDD_XCSA/X_LV1_FA1/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXADDER/Xa06/Xrb2/M4 N_XADDER/P5_XADDER/Xa06/Xrb2/M4_d
+ N_XADDER/XA06/XRB2/N002_XADDER/Xa06/Xrb2/M4_g N_VDD_XADDER/Xa06/Xrb2/M4_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA3/X_xor/M5 N_XCSA/X_LV2_HA3/X_XOR/N002_XCSA/X_LV2_HA3/X_xor/M5_d
+ N_XCSA/LV1_S[5]_XCSA/X_LV2_HA3/X_xor/M5_g
+ N_XCSA/X_LV2_HA3/X_XOR/N001_XCSA/X_LV2_HA3/X_xor/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa2/M10 N_C[3]_XCSA/Xdffa2/M10_d N_XCSA/XDFFA2/N3_XCSA/Xdffa2/M10_g
+ N_VDD_XCSA/Xdffa2/M10_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa15/M10 N_S[3]_XCSA/Xdffa15/M10_d N_XCSA/XDFFA15/N3_XCSA/Xdffa15/M10_g
+ N_VDD_XCSA/Xdffa15/M10_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel22/M6 N_XBOOTH/XSEL22/N002_XBOOTH/Xsel22/M6_d
+ N_XBOOTH/D2_XBOOTH/Xsel22/M6_g N_noxref_1594_XBOOTH/Xsel22/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel12/M6 N_XBOOTH/XSEL12/N002_XBOOTH/Xsel12/M6_d
+ N_XBOOTH/D1_XBOOTH/Xsel12/M6_g N_noxref_1595_XBOOTH/Xsel12/M6_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel02/M6 N_XBOOTH/XSEL02/N002_XBOOTH/Xsel02/M6_d
+ N_XBOOTH/D0_XBOOTH/Xsel02/M6_g N_noxref_1596_XBOOTH/Xsel02/M6_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXADDER/Xa15/Xyb3/M35 N_XADDER/XA15/XYB3/N007_XADDER/Xa15/Xyb3/M35_d
+ N_XADDER/G5_XADDER/Xa15/Xyb3/M35_g N_VDD_XADDER/Xa15/Xyb3/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXADDER/Xa64/Xao2/Xor1/M15 N_VDD_XADDER/Xa64/Xao2/Xor1/M15_d
+ N_XADDER/XA64/XAO2/N008_XADDER/Xa64/Xao2/Xor1/M15_g
+ N_XADDER/GX6[1]_XADDER/Xa64/Xao2/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mXCSA/X_LV2_HA3/M10 N_XCSA/X_LV2_HA3/N001_XCSA/X_LV2_HA3/M10_d
+ N_XCSA/LV1_S[5]_XCSA/X_LV2_HA3/M10_g N_VDD_XCSA/X_LV2_HA3/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV3_FA1/M28 N_XCSA/LV3_C[4]_XCSA/X_LV3_FA1/M28_d
+ N_XCSA/X_LV3_FA1/_COUT_XCSA/X_LV3_FA1/M28_g N_VDD_XCSA/X_LV3_FA1/M28_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXCSA/X_LV1_FA1/M4 N_XCSA/X_LV1_FA1/N001_XCSA/X_LV1_FA1/M4_d
+ N_PP1[3]_XCSA/X_LV1_FA1/M4_g N_VDD_XCSA/X_LV1_FA1/M4_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA1/M2 N_XCSA/X_LV1_FA1/_COUT_XCSA/X_LV1_FA1/M2_d
+ N_PP1[3]_XCSA/X_LV1_FA1/M2_g N_XCSA/X_LV1_FA1/P001_XCSA/X_LV1_FA1/M2_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV1_FA1/M11 N_XCSA/X_LV1_FA1/P003_XCSA/X_LV1_FA1/M11_d
+ N_PP1[3]_XCSA/X_LV1_FA1/M11_g N_XCSA/X_LV1_FA1/P002_XCSA/X_LV1_FA1/M11_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA1/M8 N_XCSA/X_LV1_FA1/N002_XCSA/X_LV1_FA1/M8_d
+ N_PP1[3]_XCSA/X_LV1_FA1/M8_g N_VDD_XCSA/X_LV1_FA1/M8_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mX02/xd27/M1 N_X02/XD27/P001_X02/xd27/M1_d N_OUT1[6]_X02/xd27/M1_g
+ N_VDD_X02/xd27/M1_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14
+ AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel22/M7 N_noxref_1594_XBOOTH/Xsel22/M7_d
+ N_XBOOTH/S2_XBOOTH/Xsel22/M7_g N_VDD_XBOOTH/Xsel22/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel12/M7 N_noxref_1595_XBOOTH/Xsel12/M7_d
+ N_XBOOTH/S1_XBOOTH/Xsel12/M7_g N_VDD_XBOOTH/Xsel12/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel02/M7 N_noxref_1596_XBOOTH/Xsel02/M7_d
+ N_XBOOTH/S0_XBOOTH/Xsel02/M7_g N_VDD_XBOOTH/Xsel02/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xdffb2/M1 N_XBOOTH/XDFFB2/P001_XBOOTH/Xdffb2/M1_d
+ N_B[2]_XBOOTH/Xdffb2/M1_g N_VDD_XBOOTH/Xdffb2/M1_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=7.7e-14 AS=2.695e-13 PD=2.8e-07 PS=1.53e-06
mXADDER/Xa15/Xyb3/Xor1/M15 N_VDD_XADDER/Xa15/Xyb3/Xor1/M15_d
+ N_XADDER/XA15/XYB3/N008_XADDER/Xa15/Xyb3/Xor1/M15_g
+ N_XADDER/GG5_XADDER/Xa15/Xyb3/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mXCSA/X_LV3_FA1/M9 N_XCSA/X_LV3_FA1/_SUM_XCSA/X_LV3_FA1/M9_d
+ N_XCSA/X_LV3_FA1/_COUT_XCSA/X_LV3_FA1/M9_g
+ N_XCSA/X_LV3_FA1/N002_XCSA/X_LV3_FA1/M9_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mX02/xd27/M2 N_X02/XD27/N0_X02/xd27/M2_d N_CLK_X02/xd27/M2_g
+ N_X02/XD27/P001_X02/xd27/M2_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV1_FA1/M5 N_XCSA/X_LV1_FA1/_COUT_XCSA/X_LV1_FA1/M5_d
+ N_PP2[1]_XCSA/X_LV1_FA1/M5_g N_XCSA/X_LV1_FA1/N001_XCSA/X_LV1_FA1/M5_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV1_FA1/M12 N_XCSA/X_LV1_FA1/_SUM_XCSA/X_LV1_FA1/M12_d
+ N_PP2[1]_XCSA/X_LV1_FA1/M12_g N_XCSA/X_LV1_FA1/P003_XCSA/X_LV1_FA1/M12_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV1_FA1/M6 N_XCSA/X_LV1_FA1/N002_XCSA/X_LV1_FA1/M6_d
+ N_PP2[1]_XCSA/X_LV1_FA1/M6_g N_VDD_XCSA/X_LV1_FA1/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXBOOTH/Xdffb2/M2 N_XBOOTH/XDFFB2/N0_XBOOTH/Xdffb2/M2_d N_CLK_XBOOTH/Xdffb2/M2_g
+ N_XBOOTH/XDFFB2/P001_XBOOTH/Xdffb2/M2_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=7.7e-14 PD=1.53e-06 PS=2.8e-07
mXCSA/Xdffa3/M1 N_XCSA/XDFFA3/P001_XCSA/Xdffa3/M1_d
+ N_XCSA/LV3_C[4]_XCSA/Xdffa3/M1_g N_VDD_XCSA/Xdffa3/M1_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa16/M1 N_XCSA/XDFFA16/P001_XCSA/Xdffa16/M1_d
+ N_XCSA/LV3_S[4]_XCSA/Xdffa16/M1_g N_VDD_XCSA/Xdffa16/M1_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXADDER/Xa37/Xao1/M11 N_XADDER/XA37/XAO1/N003_XADDER/Xa37/Xao1/M11_d
+ N_XADDER/GGG3_XADDER/Xa37/Xao1/M11_g N_VDD_XADDER/Xa37/Xao1/M11_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.474e-13
+ PD=1.42e-06 PS=6.7e-07
mXADDER/Xa06/Xrb2/M5 N_XADDER/XA06/XRB2/N001_XADDER/Xa06/Xrb2/M5_d
+ N_C[5]_XADDER/Xa06/Xrb2/M5_g N_VDD_XADDER/Xa06/Xrb2/M5_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.904e-13
+ PD=2.8e-07 PS=1.76e-06
mXBOOTH/Xsel22/M9 N_noxref_1594_XBOOTH/Xsel22/M9_d
+ N_XBOOTH/B_D[2]_XBOOTH/Xsel22/M9_g N_VDD_XBOOTH/Xsel22/M9_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel12/M9 N_noxref_1595_XBOOTH/Xsel12/M9_d
+ N_XBOOTH/B_D[2]_XBOOTH/Xsel12/M9_g N_VDD_XBOOTH/Xsel12/M9_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel02/M9 N_noxref_1596_XBOOTH/Xsel02/M9_d
+ N_XBOOTH/B_D[2]_XBOOTH/Xsel02/M9_g N_VDD_XBOOTH/Xsel02/M9_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV2_HA3/M13 N_XCSA/LV2_C[6]_XCSA/X_LV2_HA3/M13_d
+ N_XCSA/X_LV2_HA3/N001_XCSA/X_LV2_HA3/M13_g N_VDD_XCSA/X_LV2_HA3/M13_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA3/X_xor/M4 N_XCSA/LV2_S[5]_XCSA/X_LV2_HA3/X_xor/M4_d
+ N_XCSA/X_LV2_HA3/X_XOR/N002_XCSA/X_LV2_HA3/X_xor/M4_g
+ N_VDD_XCSA/X_LV2_HA3/X_xor/M4_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA1/M5 N_XCSA/X_LV3_FA1/_COUT_XCSA/X_LV3_FA1/M5_d
+ N_CACC[3]_XCSA/X_LV3_FA1/M5_g N_XCSA/X_LV3_FA1/N001_XCSA/X_LV3_FA1/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA1/M12 N_XCSA/X_LV3_FA1/_SUM_XCSA/X_LV3_FA1/M12_d
+ N_CACC[3]_XCSA/X_LV3_FA1/M12_g N_XCSA/X_LV3_FA1/P003_XCSA/X_LV3_FA1/M12_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA1/M6 N_XCSA/X_LV3_FA1/N002_XCSA/X_LV3_FA1/M6_d
+ N_CACC[3]_XCSA/X_LV3_FA1/M6_g N_VDD_XCSA/X_LV3_FA1/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/Xdffa3/M2 N_XCSA/XDFFA3/N0_XCSA/Xdffa3/M2_d N_CLK_XCSA/Xdffa3/M2_g
+ N_XCSA/XDFFA3/P001_XCSA/Xdffa3/M2_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa16/M2 N_XCSA/XDFFA16/N0_XCSA/Xdffa16/M2_d N_CLK_XCSA/Xdffa16/M2_g
+ N_XCSA/XDFFA16/P001_XCSA/Xdffa16/M2_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa06/Xrb2/M6 N_XADDER/XA06/XRB2/N002_XADDER/Xa06/Xrb2/M6_d
+ N_S[5]_XADDER/Xa06/Xrb2/M6_g N_XADDER/XA06/XRB2/N001_XADDER/Xa06/Xrb2/M6_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV1_FA1/M9 N_XCSA/X_LV1_FA1/_SUM_XCSA/X_LV1_FA1/M9_d
+ N_XCSA/X_LV1_FA1/_COUT_XCSA/X_LV1_FA1/M9_g
+ N_XCSA/X_LV1_FA1/N002_XCSA/X_LV1_FA1/M9_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXADDER/Xa27/Xyb1/Xand1/M15 N_VDD_XADDER/Xa27/Xyb1/Xand1/M15_d
+ N_XADDER/XA27/XYB1/N003_XADDER/Xa27/Xyb1/Xand1/M15_g
+ N_XADDER/PPP7_XADDER/Xa27/Xyb1/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa37/Xao1/M12 N_XADDER/XA37/XAO1/N003_XADDER/Xa37/Xao1/M12_d
+ N_XADDER/PPP7_XADDER/Xa37/Xao1/M12_g N_VDD_XADDER/Xa37/Xao1/M12_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.288e-13 AS=1.474e-13
+ PD=1.48e-06 PS=6.7e-07
mXBOOTH/Xsel22/M10 N_XBOOTH/XSEL22/B_XBOOTH/Xsel22/M10_d
+ N_XBOOTH/XSEL22/N002_XBOOTH/Xsel22/M10_g N_VDD_XBOOTH/Xsel22/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel12/M10 N_XBOOTH/XSEL12/B_XBOOTH/Xsel12/M10_d
+ N_XBOOTH/XSEL12/N002_XBOOTH/Xsel12/M10_g N_VDD_XBOOTH/Xsel12/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel02/M10 N_XBOOTH/XSEL02/B_XBOOTH/Xsel02/M10_d
+ N_XBOOTH/XSEL02/N002_XBOOTH/Xsel02/M10_g N_VDD_XBOOTH/Xsel02/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA1/M4 N_XCSA/X_LV3_FA1/N001_XCSA/X_LV3_FA1/M4_d
+ N_XCSA/LV2_S[3]_XCSA/X_LV3_FA1/M4_g N_VDD_XCSA/X_LV3_FA1/M4_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA1/M2 N_XCSA/X_LV3_FA1/_COUT_XCSA/X_LV3_FA1/M2_d
+ N_XCSA/LV2_S[3]_XCSA/X_LV3_FA1/M2_g N_XCSA/X_LV3_FA1/P001_XCSA/X_LV3_FA1/M2_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA1/M11 N_XCSA/X_LV3_FA1/P003_XCSA/X_LV3_FA1/M11_d
+ N_XCSA/LV2_S[3]_XCSA/X_LV3_FA1/M11_g
+ N_XCSA/X_LV3_FA1/P002_XCSA/X_LV3_FA1/M11_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA1/M8 N_XCSA/X_LV3_FA1/N002_XCSA/X_LV3_FA1/M8_d
+ N_XCSA/LV2_S[3]_XCSA/X_LV3_FA1/M8_g N_VDD_XCSA/X_LV3_FA1/M8_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mX02/xd27/M4 N_X02/XD27/N1_X02/xd27/M4_d N_CLK_X02/xd27/M4_g N_VDD_X02/xd27/M4_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA1/M28 N_XCSA/LV1_C[6]_XCSA/X_LV1_FA1/M28_d
+ N_XCSA/X_LV1_FA1/_COUT_XCSA/X_LV1_FA1/M28_g N_VDD_XCSA/X_LV1_FA1/M28_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXBOOTH/Xdffb2/M4 N_XBOOTH/XDFFB2/N1_XBOOTH/Xdffb2/M4_d N_CLK_XBOOTH/Xdffb2/M4_g
+ N_VDD_XBOOTH/Xdffb2/M4_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07
+ AD=2.695e-13 AS=1.485e-13 PD=1.53e-06 PS=5.4e-07
mXCSA/Xdffa3/M4 N_XCSA/XDFFA3/N1_XCSA/Xdffa3/M4_d N_CLK_XCSA/Xdffa3/M4_g
+ N_VDD_XCSA/Xdffa3/M4_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa16/M4 N_XCSA/XDFFA16/N1_XCSA/Xdffa16/M4_d N_CLK_XCSA/Xdffa16/M4_g
+ N_VDD_XCSA/Xdffa16/M4_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA1/M3 N_XCSA/X_LV3_FA1/N001_XCSA/X_LV3_FA1/M3_d
+ N_XCSA/LV2_C[3]_XCSA/X_LV3_FA1/M3_g N_VDD_XCSA/X_LV3_FA1/M3_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA1/M1 N_XCSA/X_LV3_FA1/P001_XCSA/X_LV3_FA1/M1_d
+ N_XCSA/LV2_C[3]_XCSA/X_LV3_FA1/M1_g N_VDD_XCSA/X_LV3_FA1/M1_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA1/M10 N_XCSA/X_LV3_FA1/P002_XCSA/X_LV3_FA1/M10_d
+ N_XCSA/LV2_C[3]_XCSA/X_LV3_FA1/M10_g N_VDD_XCSA/X_LV3_FA1/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA1/M7 N_XCSA/X_LV3_FA1/N002_XCSA/X_LV3_FA1/M7_d
+ N_XCSA/LV2_C[3]_XCSA/X_LV3_FA1/M7_g N_VDD_XCSA/X_LV3_FA1/M7_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mX02/xd27/M7 N_X02/XD27/N3_X02/xd27/M7_d N_X02/XD27/N1_X02/xd27/M7_g
+ N_VDD_X02/xd27/M7_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA1/M27 N_XCSA/LV1_S[5]_XCSA/X_LV1_FA1/M27_d
+ N_XCSA/X_LV1_FA1/_SUM_XCSA/X_LV1_FA1/M27_g N_VDD_XCSA/X_LV1_FA1/M27_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXBOOTH/Xdffb2/M7 N_XBOOTH/XDFFB2/N3_XBOOTH/Xdffb2/M7_d
+ N_XBOOTH/XDFFB2/N1_XBOOTH/Xdffb2/M7_g N_VDD_XBOOTH/Xdffb2/M7_s
+ N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXADDER/Xa06/Xrb1/M12 N_XADDER/XA06/XRB1/N003_XADDER/Xa06/Xrb1/M12_d
+ N_S[5]_XADDER/Xa06/Xrb1/M12_g N_VDD_XADDER/Xa06/Xrb1/M12_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa27/Xyb1/M11 N_XADDER/XA27/XYB1/N003_XADDER/Xa27/Xyb1/M11_d
+ N_XADDER/PP5_XADDER/Xa27/Xyb1/M11_g N_VDD_XADDER/Xa27/Xyb1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mXADDER/Xa37/Xao1/Xand1/M15 N_VDD_XADDER/Xa37/Xao1/Xand1/M15_d
+ N_XADDER/XA37/XAO1/N003_XADDER/Xa37/Xao1/Xand1/M15_g
+ N_XADDER/XA37/OUT1_XADDER/Xa37/Xao1/Xand1/M15_s N_VDD_XADDER/Xa72/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa3/M7 N_XCSA/XDFFA3/N3_XCSA/Xdffa3/M7_d
+ N_XCSA/XDFFA3/N1_XCSA/Xdffa3/M7_g N_VDD_XCSA/Xdffa3/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa16/M7 N_XCSA/XDFFA16/N3_XCSA/Xdffa16/M7_d
+ N_XCSA/XDFFA16/N1_XCSA/Xdffa16/M7_g N_VDD_XCSA/Xdffa16/M7_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel22/M16 N_XBOOTH/XSEL22/N003_XBOOTH/Xsel22/M16_d
+ N_A_D[5]_XBOOTH/Xsel22/M16_g N_VDD_XBOOTH/Xsel22/M16_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel12/M16 N_XBOOTH/XSEL12/N003_XBOOTH/Xsel12/M16_d
+ N_A_D[3]_XBOOTH/Xsel12/M16_g N_VDD_XBOOTH/Xsel12/M16_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel02/M16 N_XBOOTH/XSEL02/N003_XBOOTH/Xsel02/M16_d
+ N_A_D[1]_XBOOTH/Xsel02/M16_g N_VDD_XBOOTH/Xsel02/M16_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXADDER/Xa06/Xrb1/M11 N_XADDER/XA06/XRB1/N003_XADDER/Xa06/Xrb1/M11_d
+ N_C[5]_XADDER/Xa06/Xrb1/M11_g N_VDD_XADDER/Xa06/Xrb1/M11_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa27/Xyb1/M12 N_XADDER/XA27/XYB1/N003_XADDER/Xa27/Xyb1/M12_d
+ N_XADDER/PP7_XADDER/Xa27/Xyb1/M12_g N_VDD_XADDER/Xa27/Xyb1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel22/M15 N_XBOOTH/XSEL22/N004_XBOOTH/Xsel22/M15_d
+ N_XBOOTH/XSEL22/B_XBOOTH/Xsel22/M15_g N_XBOOTH/XSEL22/N003_XBOOTH/Xsel22/M15_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel12/M15 N_XBOOTH/XSEL12/N004_XBOOTH/Xsel12/M15_d
+ N_XBOOTH/XSEL12/B_XBOOTH/Xsel12/M15_g N_XBOOTH/XSEL12/N003_XBOOTH/Xsel12/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel02/M15 N_XBOOTH/XSEL02/N004_XBOOTH/Xsel02/M15_d
+ N_XBOOTH/XSEL02/B_XBOOTH/Xsel02/M15_g N_XBOOTH/XSEL02/N003_XBOOTH/Xsel02/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mX02/xd27/M10 N_OUT[6]_X02/xd27/M10_d N_X02/XD27/N3_X02/xd27/M10_g
+ N_VDD_X02/xd27/M10_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA2/M27 N_XCSA/LV3_S[4]_XCSA/X_LV3_FA2/M27_d
+ N_XCSA/X_LV3_FA2/_SUM_XCSA/X_LV3_FA2/M27_g N_VDD_XCSA/X_LV3_FA2/M27_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXBOOTH/Xdffb2/M10 N_XBOOTH/B_D[2]_XBOOTH/Xdffb2/M10_d
+ N_XBOOTH/XDFFB2/N3_XBOOTH/Xdffb2/M10_g N_VDD_XBOOTH/Xdffb2/M10_s
+ N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa37/Xao2/M36 N_XADDER/XA37/XAO2/N008_XADDER/Xa37/Xao2/M36_d
+ N_XADDER/XA37/OUT1_XADDER/Xa37/Xao2/M36_g
+ N_XADDER/XA37/XAO2/N007_XADDER/Xa37/Xao2/M36_s N_VDD_XADDER/Xa72/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXCSA/Xdffa3/M10 N_C[4]_XCSA/Xdffa3/M10_d N_XCSA/XDFFA3/N3_XCSA/Xdffa3/M10_g
+ N_VDD_XCSA/Xdffa3/M10_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa16/M10 N_S[4]_XCSA/Xdffa16/M10_d N_XCSA/XDFFA16/N3_XCSA/Xdffa16/M10_g
+ N_VDD_XCSA/Xdffa16/M10_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA4/M9 N_XCSA/X_LV2_HA4/N001_XCSA/X_LV2_HA4/M9_d
+ N_XCSA/LV1_C[6]_XCSA/X_LV2_HA4/M9_g N_VDD_XCSA/X_LV2_HA4/M9_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA4/X_xor/M6 N_XCSA/X_LV2_HA4/X_XOR/N001_XCSA/X_LV2_HA4/X_xor/M6_d
+ N_XCSA/LV1_C[6]_XCSA/X_LV2_HA4/X_xor/M6_g N_VDD_XCSA/X_LV2_HA4/X_xor/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV1_FA2/M3 N_XCSA/X_LV1_FA2/N001_XCSA/X_LV1_FA2/M3_d
+ N_PP0[6]_XCSA/X_LV1_FA2/M3_g N_VDD_XCSA/X_LV1_FA2/M3_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV1_FA2/M1 N_XCSA/X_LV1_FA2/P001_XCSA/X_LV1_FA2/M1_d
+ N_PP0[6]_XCSA/X_LV1_FA2/M1_g N_VDD_XCSA/X_LV1_FA2/M1_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV1_FA2/M10 N_XCSA/X_LV1_FA2/P002_XCSA/X_LV1_FA2/M10_d
+ N_PP0[6]_XCSA/X_LV1_FA2/M10_g N_VDD_XCSA/X_LV1_FA2/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV1_FA2/M7 N_XCSA/X_LV1_FA2/N002_XCSA/X_LV1_FA2/M7_d
+ N_PP0[6]_XCSA/X_LV1_FA2/M7_g N_VDD_XCSA/X_LV1_FA2/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA2/M28 N_XCSA/LV3_C[5]_XCSA/X_LV3_FA2/M28_d
+ N_XCSA/X_LV3_FA2/_COUT_XCSA/X_LV3_FA2/M28_g N_VDD_XCSA/X_LV3_FA2/M28_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa06/Xrb1/Xand1/M15 N_VDD_XADDER/Xa06/Xrb1/Xand1/M15_d
+ N_XADDER/XA06/XRB1/N003_XADDER/Xa06/Xrb1/Xand1/M15_g
+ N_XADDER/G5_XADDER/Xa06/Xrb1/Xand1/M15_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa27/Xyb2/M12 N_XADDER/XA27/XYB2/N003_XADDER/Xa27/Xyb2/M12_d
+ N_XADDER/PP7_XADDER/Xa27/Xyb2/M12_g N_VDD_XADDER/Xa27/Xyb2/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa37/Xao2/M35 N_XADDER/XA37/XAO2/N007_XADDER/Xa37/Xao2/M35_d
+ N_XADDER/GGG7_XADDER/Xa37/Xao2/M35_g N_VDD_XADDER/Xa37/Xao2/M35_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXBOOTH/Xsel22/M14 N_PP2[2]_XBOOTH/Xsel22/M14_d
+ N_XBOOTH/XSEL22/N004_XBOOTH/Xsel22/M14_g N_VDD_XBOOTH/Xsel22/M14_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel12/M14 N_PP1[2]_XBOOTH/Xsel12/M14_d
+ N_XBOOTH/XSEL12/N004_XBOOTH/Xsel12/M14_g N_VDD_XBOOTH/Xsel12/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel02/M14 N_PP0[2]_XBOOTH/Xsel02/M14_d
+ N_XBOOTH/XSEL02/N004_XBOOTH/Xsel02/M14_g N_VDD_XBOOTH/Xsel02/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA4/X_xor/M5 N_XCSA/X_LV2_HA4/X_XOR/N002_XCSA/X_LV2_HA4/X_xor/M5_d
+ N_XCSA/LV1_S[6]_XCSA/X_LV2_HA4/X_xor/M5_g
+ N_XCSA/X_LV2_HA4/X_XOR/N001_XCSA/X_LV2_HA4/X_xor/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV3_FA2/M9 N_XCSA/X_LV3_FA2/_SUM_XCSA/X_LV3_FA2/M9_d
+ N_XCSA/X_LV3_FA2/_COUT_XCSA/X_LV3_FA2/M9_g
+ N_XCSA/X_LV3_FA2/N002_XCSA/X_LV3_FA2/M9_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXCSA/X_LV2_HA4/M10 N_XCSA/X_LV2_HA4/N001_XCSA/X_LV2_HA4/M10_d
+ N_XCSA/LV1_S[6]_XCSA/X_LV2_HA4/M10_g N_VDD_XCSA/X_LV2_HA4/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA2/M4 N_XCSA/X_LV1_FA2/N001_XCSA/X_LV1_FA2/M4_d
+ N_PP1[4]_XCSA/X_LV1_FA2/M4_g N_VDD_XCSA/X_LV1_FA2/M4_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA2/M2 N_XCSA/X_LV1_FA2/_COUT_XCSA/X_LV1_FA2/M2_d
+ N_PP1[4]_XCSA/X_LV1_FA2/M2_g N_XCSA/X_LV1_FA2/P001_XCSA/X_LV1_FA2/M2_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV1_FA2/M11 N_XCSA/X_LV1_FA2/P003_XCSA/X_LV1_FA2/M11_d
+ N_PP1[4]_XCSA/X_LV1_FA2/M11_g N_XCSA/X_LV1_FA2/P002_XCSA/X_LV1_FA2/M11_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA2/M8 N_XCSA/X_LV1_FA2/N002_XCSA/X_LV1_FA2/M8_d
+ N_PP1[4]_XCSA/X_LV1_FA2/M8_g N_VDD_XCSA/X_LV1_FA2/M8_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mXADDER/Xa27/Xyb2/M11 N_XADDER/XA27/XYB2/N003_XADDER/Xa27/Xyb2/M11_d
+ N_XADDER/GG5_XADDER/Xa27/Xyb2/M11_g N_VDD_XADDER/Xa27/Xyb2/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mXADDER/Xa37/Xao2/Xor1/M15 N_VDD_XADDER/Xa37/Xao2/Xor1/M15_d
+ N_XADDER/XA37/XAO2/N008_XADDER/Xa37/Xao2/Xor1/M15_g
+ N_XADDER/GOUT7_XADDER/Xa37/Xao2/Xor1/M15_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mXCSA/Xdffa4/M1 N_XCSA/XDFFA4/P001_XCSA/Xdffa4/M1_d
+ N_XCSA/LV3_C[5]_XCSA/Xdffa4/M1_g N_VDD_XCSA/Xdffa4/M1_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa17/M1 N_XCSA/XDFFA17/P001_XCSA/Xdffa17/M1_d
+ N_XCSA/LV3_S[5]_XCSA/Xdffa17/M1_g N_VDD_XCSA/Xdffa17/M1_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXADDER/Xa17/Xyb1/Xand1/M15 N_VDD_XADDER/Xa17/Xyb1/Xand1/M15_d
+ N_XADDER/XA17/XYB1/N003_XADDER/Xa17/Xyb1/Xand1/M15_g
+ N_XADDER/PP7_XADDER/Xa17/Xyb1/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA2/M5 N_XCSA/X_LV1_FA2/_COUT_XCSA/X_LV1_FA2/M5_d
+ N_PP2[2]_XCSA/X_LV1_FA2/M5_g N_XCSA/X_LV1_FA2/N001_XCSA/X_LV1_FA2/M5_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV1_FA2/M12 N_XCSA/X_LV1_FA2/_SUM_XCSA/X_LV1_FA2/M12_d
+ N_PP2[2]_XCSA/X_LV1_FA2/M12_g N_XCSA/X_LV1_FA2/P003_XCSA/X_LV1_FA2/M12_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV1_FA2/M6 N_XCSA/X_LV1_FA2/N002_XCSA/X_LV1_FA2/M6_d
+ N_PP2[2]_XCSA/X_LV1_FA2/M6_g N_VDD_XCSA/X_LV1_FA2/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA2/M5 N_XCSA/X_LV3_FA2/_COUT_XCSA/X_LV3_FA2/M5_d
+ N_CACC[4]_XCSA/X_LV3_FA2/M5_g N_XCSA/X_LV3_FA2/N001_XCSA/X_LV3_FA2/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA2/M12 N_XCSA/X_LV3_FA2/_SUM_XCSA/X_LV3_FA2/M12_d
+ N_CACC[4]_XCSA/X_LV3_FA2/M12_g N_XCSA/X_LV3_FA2/P003_XCSA/X_LV3_FA2/M12_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA2/M6 N_XCSA/X_LV3_FA2/N002_XCSA/X_LV3_FA2/M6_d
+ N_CACC[4]_XCSA/X_LV3_FA2/M6_g N_VDD_XCSA/X_LV3_FA2/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXADDER/Xa07/Xrb2/M4 N_XADDER/P6_XADDER/Xa07/Xrb2/M4_d
+ N_XADDER/XA07/XRB2/N002_XADDER/Xa07/Xrb2/M4_g N_VDD_XADDER/Xa07/Xrb2/M4_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa4/M2 N_XCSA/XDFFA4/N0_XCSA/Xdffa4/M2_d N_CLK_XCSA/Xdffa4/M2_g
+ N_XCSA/XDFFA4/P001_XCSA/Xdffa4/M2_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa17/M2 N_XCSA/XDFFA17/N0_XCSA/Xdffa17/M2_d N_CLK_XCSA/Xdffa17/M2_g
+ N_XCSA/XDFFA17/P001_XCSA/Xdffa17/M2_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV2_HA4/M13 N_XCSA/LV2_C[7]_XCSA/X_LV2_HA4/M13_d
+ N_XCSA/X_LV2_HA4/N001_XCSA/X_LV2_HA4/M13_g N_VDD_XCSA/X_LV2_HA4/M13_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA4/X_xor/M4 N_XCSA/LV2_S[6]_XCSA/X_LV2_HA4/X_xor/M4_d
+ N_XCSA/X_LV2_HA4/X_XOR/N002_XCSA/X_LV2_HA4/X_xor/M4_g
+ N_VDD_XCSA/X_LV2_HA4/X_xor/M4_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA2/M4 N_XCSA/X_LV3_FA2/N001_XCSA/X_LV3_FA2/M4_d
+ N_XCSA/LV2_S[4]_XCSA/X_LV3_FA2/M4_g N_VDD_XCSA/X_LV3_FA2/M4_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA2/M2 N_XCSA/X_LV3_FA2/_COUT_XCSA/X_LV3_FA2/M2_d
+ N_XCSA/LV2_S[4]_XCSA/X_LV3_FA2/M2_g N_XCSA/X_LV3_FA2/P001_XCSA/X_LV3_FA2/M2_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA2/M11 N_XCSA/X_LV3_FA2/P003_XCSA/X_LV3_FA2/M11_d
+ N_XCSA/LV2_S[4]_XCSA/X_LV3_FA2/M11_g
+ N_XCSA/X_LV3_FA2/P002_XCSA/X_LV3_FA2/M11_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA2/M8 N_XCSA/X_LV3_FA2/N002_XCSA/X_LV3_FA2/M8_d
+ N_XCSA/LV2_S[4]_XCSA/X_LV3_FA2/M8_g N_VDD_XCSA/X_LV3_FA2/M8_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV1_FA2/M9 N_XCSA/X_LV1_FA2/_SUM_XCSA/X_LV1_FA2/M9_d
+ N_XCSA/X_LV1_FA2/_COUT_XCSA/X_LV1_FA2/M9_g
+ N_XCSA/X_LV1_FA2/N002_XCSA/X_LV1_FA2/M9_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXADDER/Xa27/Xyb2/Xand1/M15 N_VDD_XADDER/Xa27/Xyb2/Xand1/M15_d
+ N_XADDER/XA27/XYB2/N003_XADDER/Xa27/Xyb2/Xand1/M15_g
+ N_XADDER/XA27/T1_XADDER/Xa27/Xyb2/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel23/M8 N_XBOOTH/XSEL23/N002_XBOOTH/Xsel23/M8_d
+ N_XBOOTH/B_D[2]_XBOOTH/Xsel23/M8_g N_noxref_1639_XBOOTH/Xsel23/M8_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel13/M8 N_XBOOTH/XSEL13/N002_XBOOTH/Xsel13/M8_d
+ N_XBOOTH/B_D[2]_XBOOTH/Xsel13/M8_g N_noxref_1640_XBOOTH/Xsel13/M8_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel03/M8 N_XBOOTH/XSEL03/N002_XBOOTH/Xsel03/M8_d
+ N_XBOOTH/B_D[2]_XBOOTH/Xsel03/M8_g N_noxref_1641_XBOOTH/Xsel03/M8_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_FA2/M28 N_XCSA/LV1_C[7]_XCSA/X_LV1_FA2/M28_d
+ N_XCSA/X_LV1_FA2/_COUT_XCSA/X_LV1_FA2/M28_g N_VDD_XCSA/X_LV1_FA2/M28_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa17/Xyb1/M11 N_XADDER/XA17/XYB1/N003_XADDER/Xa17/Xyb1/M11_d
+ N_XADDER/P6_XADDER/Xa17/Xyb1/M11_g N_VDD_XADDER/Xa17/Xyb1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mXCSA/X_LV3_FA2/M3 N_XCSA/X_LV3_FA2/N001_XCSA/X_LV3_FA2/M3_d
+ N_XCSA/LV2_C[4]_XCSA/X_LV3_FA2/M3_g N_VDD_XCSA/X_LV3_FA2/M3_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA2/M1 N_XCSA/X_LV3_FA2/P001_XCSA/X_LV3_FA2/M1_d
+ N_XCSA/LV2_C[4]_XCSA/X_LV3_FA2/M1_g N_VDD_XCSA/X_LV3_FA2/M1_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA2/M10 N_XCSA/X_LV3_FA2/P002_XCSA/X_LV3_FA2/M10_d
+ N_XCSA/LV2_C[4]_XCSA/X_LV3_FA2/M10_g N_VDD_XCSA/X_LV3_FA2/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA2/M7 N_XCSA/X_LV3_FA2/N002_XCSA/X_LV3_FA2/M7_d
+ N_XCSA/LV2_C[4]_XCSA/X_LV3_FA2/M7_g N_VDD_XCSA/X_LV3_FA2/M7_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/Xdffa4/M4 N_XCSA/XDFFA4/N1_XCSA/Xdffa4/M4_d N_CLK_XCSA/Xdffa4/M4_g
+ N_VDD_XCSA/Xdffa4/M4_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa17/M4 N_XCSA/XDFFA17/N1_XCSA/Xdffa17/M4_d N_CLK_XCSA/Xdffa17/M4_g
+ N_VDD_XCSA/Xdffa17/M4_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXADDER/Xa07/Xrb2/M5 N_XADDER/XA07/XRB2/N001_XADDER/Xa07/Xrb2/M5_d
+ N_C[6]_XADDER/Xa07/Xrb2/M5_g N_VDD_XADDER/Xa07/Xrb2/M5_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.904e-13
+ PD=2.8e-07 PS=1.76e-06
mXBOOTH/Xsel23/M6 N_XBOOTH/XSEL23/N002_XBOOTH/Xsel23/M6_d
+ N_XBOOTH/D2_XBOOTH/Xsel23/M6_g N_noxref_1639_XBOOTH/Xsel23/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel13/M6 N_XBOOTH/XSEL13/N002_XBOOTH/Xsel13/M6_d
+ N_XBOOTH/D1_XBOOTH/Xsel13/M6_g N_noxref_1640_XBOOTH/Xsel13/M6_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel03/M6 N_XBOOTH/XSEL03/N002_XBOOTH/Xsel03/M6_d
+ N_XBOOTH/D0_XBOOTH/Xsel03/M6_g N_noxref_1641_XBOOTH/Xsel03/M6_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXADDER/Xa17/Xyb1/M12 N_XADDER/XA17/XYB1/N003_XADDER/Xa17/Xyb1/M12_d
+ N_XADDER/P7_XADDER/Xa17/Xyb1/M12_g N_VDD_XADDER/Xa17/Xyb1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA2/M27 N_XCSA/LV1_S[6]_XCSA/X_LV1_FA2/M27_d
+ N_XCSA/X_LV1_FA2/_SUM_XCSA/X_LV1_FA2/M27_g N_VDD_XCSA/X_LV1_FA2/M27_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXBOOTH/Xdffb3/M1 N_XBOOTH/XDFFB3/P001_XBOOTH/Xdffb3/M1_d
+ N_B[3]_XBOOTH/Xdffb3/M1_g N_VDD_XBOOTH/Xdffb3/M1_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=7.7e-14 AS=2.695e-13 PD=2.8e-07 PS=1.53e-06
mXADDER/Xa07/Xrb2/M6 N_XADDER/XA07/XRB2/N002_XADDER/Xa07/Xrb2/M6_d
+ N_S[6]_XADDER/Xa07/Xrb2/M6_g N_XADDER/XA07/XRB2/N001_XADDER/Xa07/Xrb2/M6_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa4/M7 N_XCSA/XDFFA4/N3_XCSA/Xdffa4/M7_d
+ N_XCSA/XDFFA4/N1_XCSA/Xdffa4/M7_g N_VDD_XCSA/Xdffa4/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa17/M7 N_XCSA/XDFFA17/N3_XCSA/Xdffa17/M7_d
+ N_XCSA/XDFFA17/N1_XCSA/Xdffa17/M7_g N_VDD_XCSA/Xdffa17/M7_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa27/Xyb3/M36 N_XADDER/XA27/XYB3/N008_XADDER/Xa27/Xyb3/M36_d
+ N_XADDER/XA27/T1_XADDER/Xa27/Xyb3/M36_g
+ N_XADDER/XA27/XYB3/N007_XADDER/Xa27/Xyb3/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXBOOTH/Xsel23/M7 N_noxref_1639_XBOOTH/Xsel23/M7_d
+ N_XBOOTH/S2_XBOOTH/Xsel23/M7_g N_VDD_XBOOTH/Xsel23/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel13/M7 N_noxref_1640_XBOOTH/Xsel13/M7_d
+ N_XBOOTH/S1_XBOOTH/Xsel13/M7_g N_VDD_XBOOTH/Xsel13/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel03/M7 N_noxref_1641_XBOOTH/Xsel03/M7_d
+ N_XBOOTH/S0_XBOOTH/Xsel03/M7_g N_VDD_XBOOTH/Xsel03/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xdffb3/M2 N_XBOOTH/XDFFB3/N0_XBOOTH/Xdffb3/M2_d N_CLK_XBOOTH/Xdffb3/M2_g
+ N_XBOOTH/XDFFB3/P001_XBOOTH/Xdffb3/M2_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=7.7e-14 PD=1.53e-06 PS=2.8e-07
mXCSA/X_LV3_FA3/M27 N_XCSA/LV3_S[5]_XCSA/X_LV3_FA3/M27_d
+ N_XCSA/X_LV3_FA3/_SUM_XCSA/X_LV3_FA3/M27_g N_VDD_XCSA/X_LV3_FA3/M27_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa27/Xyb3/M35 N_XADDER/XA27/XYB3/N007_XADDER/Xa27/Xyb3/M35_d
+ N_XADDER/GG7_XADDER/Xa27/Xyb3/M35_g N_VDD_XADDER/Xa27/Xyb3/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXBOOTH/Xsel23/M9 N_noxref_1639_XBOOTH/Xsel23/M9_d
+ N_XBOOTH/B_D[3]_XBOOTH/Xsel23/M9_g N_VDD_XBOOTH/Xsel23/M9_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel13/M9 N_noxref_1640_XBOOTH/Xsel13/M9_d
+ N_XBOOTH/B_D[3]_XBOOTH/Xsel13/M9_g N_VDD_XBOOTH/Xsel13/M9_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel03/M9 N_noxref_1641_XBOOTH/Xsel03/M9_d
+ N_XBOOTH/B_D[3]_XBOOTH/Xsel03/M9_g N_VDD_XBOOTH/Xsel03/M9_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa17/Xyb2/M12 N_XADDER/XA17/XYB2/N003_XADDER/Xa17/Xyb2/M12_d
+ N_XADDER/P7_XADDER/Xa17/Xyb2/M12_g N_VDD_XADDER/Xa17/Xyb2/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA3/M28 N_XCSA/LV3_C[6]_XCSA/X_LV3_FA3/M28_d
+ N_XCSA/X_LV3_FA3/_COUT_XCSA/X_LV3_FA3/M28_g N_VDD_XCSA/X_LV3_FA3/M28_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa07/Xrb1/M12 N_XADDER/XA07/XRB1/N003_XADDER/Xa07/Xrb1/M12_d
+ N_S[6]_XADDER/Xa07/Xrb1/M12_g N_VDD_XADDER/Xa07/Xrb1/M12_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa4/M10 N_C[5]_XCSA/Xdffa4/M10_d N_XCSA/XDFFA4/N3_XCSA/Xdffa4/M10_g
+ N_VDD_XCSA/Xdffa4/M10_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa17/M10 N_S[5]_XCSA/Xdffa17/M10_d N_XCSA/XDFFA17/N3_XCSA/Xdffa17/M10_g
+ N_VDD_XCSA/Xdffa17/M10_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa27/Xyb3/Xor1/M15 N_VDD_XADDER/Xa27/Xyb3/Xor1/M15_d
+ N_XADDER/XA27/XYB3/N008_XADDER/Xa27/Xyb3/Xor1/M15_g
+ N_XADDER/GGG7_XADDER/Xa27/Xyb3/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mXBOOTH/Xdffb3/M4 N_XBOOTH/XDFFB3/N1_XBOOTH/Xdffb3/M4_d N_CLK_XBOOTH/Xdffb3/M4_g
+ N_VDD_XBOOTH/Xdffb3/M4_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07
+ AD=2.695e-13 AS=1.485e-13 PD=1.53e-06 PS=5.4e-07
mXBOOTH/Xsel23/M10 N_XBOOTH/XSEL23/B_XBOOTH/Xsel23/M10_d
+ N_XBOOTH/XSEL23/N002_XBOOTH/Xsel23/M10_g N_VDD_XBOOTH/Xsel23/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel13/M10 N_XBOOTH/XSEL13/B_XBOOTH/Xsel13/M10_d
+ N_XBOOTH/XSEL13/N002_XBOOTH/Xsel13/M10_g N_VDD_XBOOTH/Xsel13/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel03/M10 N_XBOOTH/XSEL03/B_XBOOTH/Xsel03/M10_d
+ N_XBOOTH/XSEL03/N002_XBOOTH/Xsel03/M10_g N_VDD_XBOOTH/Xsel03/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa17/Xyb2/M11 N_XADDER/XA17/XYB2/N003_XADDER/Xa17/Xyb2/M11_d
+ N_XADDER/G6_XADDER/Xa17/Xyb2/M11_g N_VDD_XADDER/Xa17/Xyb2/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mXCSA/X_LV3_FA3/M9 N_XCSA/X_LV3_FA3/_SUM_XCSA/X_LV3_FA3/M9_d
+ N_XCSA/X_LV3_FA3/_COUT_XCSA/X_LV3_FA3/M9_g
+ N_XCSA/X_LV3_FA3/N002_XCSA/X_LV3_FA3/M9_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXCSA/X_LV1_FA3/M3 N_XCSA/X_LV1_FA3/N001_XCSA/X_LV1_FA3/M3_d
+ N_PP0[6]_XCSA/X_LV1_FA3/M3_g N_VDD_XCSA/X_LV1_FA3/M3_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV1_FA3/M1 N_XCSA/X_LV1_FA3/P001_XCSA/X_LV1_FA3/M1_d
+ N_PP0[6]_XCSA/X_LV1_FA3/M1_g N_VDD_XCSA/X_LV1_FA3/M1_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV1_FA3/M10 N_XCSA/X_LV1_FA3/P002_XCSA/X_LV1_FA3/M10_d
+ N_PP0[6]_XCSA/X_LV1_FA3/M10_g N_VDD_XCSA/X_LV1_FA3/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV1_FA3/M7 N_XCSA/X_LV1_FA3/N002_XCSA/X_LV1_FA3/M7_d
+ N_PP0[6]_XCSA/X_LV1_FA3/M7_g N_VDD_XCSA/X_LV1_FA3/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXADDER/Xa07/Xrb1/M11 N_XADDER/XA07/XRB1/N003_XADDER/Xa07/Xrb1/M11_d
+ N_C[6]_XADDER/Xa07/Xrb1/M11_g N_VDD_XADDER/Xa07/Xrb1/M11_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa76/M4 N_OUT1[6]_XADDER/Xa76/M4_d N_XADDER/XA76/N002_XADDER/Xa76/M4_g
+ N_VDD_XADDER/Xa76/M4_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd29/M1 N_X02/XD29/P001_X02/xd29/M1_d N_OUT1[8]_X02/xd29/M1_g
+ N_VDD_X02/xd29/M1_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14
+ AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xdffb3/M7 N_XBOOTH/XDFFB3/N3_XBOOTH/Xdffb3/M7_d
+ N_XBOOTH/XDFFB3/N1_XBOOTH/Xdffb3/M7_g N_VDD_XBOOTH/Xdffb3/M7_s
+ N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV2_HA5/M9 N_XCSA/X_LV2_HA5/N001_XCSA/X_LV2_HA5/M9_d
+ N_XCSA/LV1_C[7]_XCSA/X_LV2_HA5/M9_g N_VDD_XCSA/X_LV2_HA5/M9_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA5/X_xor/M6 N_XCSA/X_LV2_HA5/X_XOR/N001_XCSA/X_LV2_HA5/X_xor/M6_d
+ N_XCSA/LV1_C[7]_XCSA/X_LV2_HA5/X_xor/M6_g N_VDD_XCSA/X_LV2_HA5/X_xor/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mX02/xd29/M2 N_X02/XD29/N0_X02/xd29/M2_d N_CLK_X02/xd29/M2_g
+ N_X02/XD29/P001_X02/xd29/M2_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV1_FA3/M4 N_XCSA/X_LV1_FA3/N001_XCSA/X_LV1_FA3/M4_d
+ N_PP1[5]_XCSA/X_LV1_FA3/M4_g N_VDD_XCSA/X_LV1_FA3/M4_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA3/M2 N_XCSA/X_LV1_FA3/_COUT_XCSA/X_LV1_FA3/M2_d
+ N_PP1[5]_XCSA/X_LV1_FA3/M2_g N_XCSA/X_LV1_FA3/P001_XCSA/X_LV1_FA3/M2_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV1_FA3/M11 N_XCSA/X_LV1_FA3/P003_XCSA/X_LV1_FA3/M11_d
+ N_PP1[5]_XCSA/X_LV1_FA3/M11_g N_XCSA/X_LV1_FA3/P002_XCSA/X_LV1_FA3/M11_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA3/M8 N_XCSA/X_LV1_FA3/N002_XCSA/X_LV1_FA3/M8_d
+ N_PP1[5]_XCSA/X_LV1_FA3/M8_g N_VDD_XCSA/X_LV1_FA3/M8_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA3/M5 N_XCSA/X_LV3_FA3/_COUT_XCSA/X_LV3_FA3/M5_d
+ N_CACC[5]_XCSA/X_LV3_FA3/M5_g N_XCSA/X_LV3_FA3/N001_XCSA/X_LV3_FA3/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA3/M12 N_XCSA/X_LV3_FA3/_SUM_XCSA/X_LV3_FA3/M12_d
+ N_CACC[5]_XCSA/X_LV3_FA3/M12_g N_XCSA/X_LV3_FA3/P003_XCSA/X_LV3_FA3/M12_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA3/M6 N_XCSA/X_LV3_FA3/N002_XCSA/X_LV3_FA3/M6_d
+ N_CACC[5]_XCSA/X_LV3_FA3/M6_g N_VDD_XCSA/X_LV3_FA3/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/Xdffa5/M1 N_XCSA/XDFFA5/P001_XCSA/Xdffa5/M1_d
+ N_XCSA/LV3_C[6]_XCSA/Xdffa5/M1_g N_VDD_XCSA/Xdffa5/M1_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa18/M1 N_XCSA/XDFFA18/P001_XCSA/Xdffa18/M1_d
+ N_XCSA/LV3_S[6]_XCSA/Xdffa18/M1_g N_VDD_XCSA/Xdffa18/M1_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV2_HA5/X_xor/M5 N_XCSA/X_LV2_HA5/X_XOR/N002_XCSA/X_LV2_HA5/X_xor/M5_d
+ N_XCSA/LV1_S[7]_XCSA/X_LV2_HA5/X_xor/M5_g
+ N_XCSA/X_LV2_HA5/X_XOR/N001_XCSA/X_LV2_HA5/X_xor/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV2_HA5/M10 N_XCSA/X_LV2_HA5/N001_XCSA/X_LV2_HA5/M10_d
+ N_XCSA/LV1_S[7]_XCSA/X_LV2_HA5/M10_g N_VDD_XCSA/X_LV2_HA5/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/Xdffa5/M2 N_XCSA/XDFFA5/N0_XCSA/Xdffa5/M2_d N_CLK_XCSA/Xdffa5/M2_g
+ N_XCSA/XDFFA5/P001_XCSA/Xdffa5/M2_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa18/M2 N_XCSA/XDFFA18/N0_XCSA/Xdffa18/M2_d N_CLK_XCSA/Xdffa18/M2_g
+ N_XCSA/XDFFA18/P001_XCSA/Xdffa18/M2_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV1_FA3/M5 N_XCSA/X_LV1_FA3/_COUT_XCSA/X_LV1_FA3/M5_d
+ N_PP2[3]_XCSA/X_LV1_FA3/M5_g N_XCSA/X_LV1_FA3/N001_XCSA/X_LV1_FA3/M5_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV1_FA3/M12 N_XCSA/X_LV1_FA3/_SUM_XCSA/X_LV1_FA3/M12_d
+ N_PP2[3]_XCSA/X_LV1_FA3/M12_g N_XCSA/X_LV1_FA3/P003_XCSA/X_LV1_FA3/M12_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV1_FA3/M6 N_XCSA/X_LV1_FA3/N002_XCSA/X_LV1_FA3/M6_d
+ N_PP2[3]_XCSA/X_LV1_FA3/M6_g N_VDD_XCSA/X_LV1_FA3/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXADDER/Xa17/Xyb2/Xand1/M15 N_VDD_XADDER/Xa17/Xyb2/Xand1/M15_d
+ N_XADDER/XA17/XYB2/N003_XADDER/Xa17/Xyb2/Xand1/M15_g
+ N_XADDER/XA17/T1_XADDER/Xa17/Xyb2/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA3/M4 N_XCSA/X_LV3_FA3/N001_XCSA/X_LV3_FA3/M4_d
+ N_XCSA/LV2_S[5]_XCSA/X_LV3_FA3/M4_g N_VDD_XCSA/X_LV3_FA3/M4_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA3/M2 N_XCSA/X_LV3_FA3/_COUT_XCSA/X_LV3_FA3/M2_d
+ N_XCSA/LV2_S[5]_XCSA/X_LV3_FA3/M2_g N_XCSA/X_LV3_FA3/P001_XCSA/X_LV3_FA3/M2_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA3/M11 N_XCSA/X_LV3_FA3/P003_XCSA/X_LV3_FA3/M11_d
+ N_XCSA/LV2_S[5]_XCSA/X_LV3_FA3/M11_g
+ N_XCSA/X_LV3_FA3/P002_XCSA/X_LV3_FA3/M11_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA3/M8 N_XCSA/X_LV3_FA3/N002_XCSA/X_LV3_FA3/M8_d
+ N_XCSA/LV2_S[5]_XCSA/X_LV3_FA3/M8_g N_VDD_XCSA/X_LV3_FA3/M8_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mXBOOTH/Xsel23/M16 N_XBOOTH/XSEL23/N003_XBOOTH/Xsel23/M16_d
+ N_A_D[5]_XBOOTH/Xsel23/M16_g N_VDD_XBOOTH/Xsel23/M16_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel13/M16 N_XBOOTH/XSEL13/N003_XBOOTH/Xsel13/M16_d
+ N_A_D[3]_XBOOTH/Xsel13/M16_g N_VDD_XBOOTH/Xsel13/M16_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel03/M16 N_XBOOTH/XSEL03/N003_XBOOTH/Xsel03/M16_d
+ N_A_D[1]_XBOOTH/Xsel03/M16_g N_VDD_XBOOTH/Xsel03/M16_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXADDER/Xa07/Xrb1/Xand1/M15 N_VDD_XADDER/Xa07/Xrb1/Xand1/M15_d
+ N_XADDER/XA07/XRB1/N003_XADDER/Xa07/Xrb1/Xand1/M15_g
+ N_XADDER/G6_XADDER/Xa07/Xrb1/Xand1/M15_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa66/Xao1/M11 N_XADDER/XA66/XAO1/N003_XADDER/Xa66/Xao1/M11_d
+ N_XADDER/GX5[0]_XADDER/Xa66/Xao1/M11_g N_VDD_XADDER/Xa66/Xao1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.474e-13
+ PD=1.42e-06 PS=6.7e-07
mXBOOTH/Xdffb3/M10 N_XBOOTH/B_D[3]_XBOOTH/Xdffb3/M10_d
+ N_XBOOTH/XDFFB3/N3_XBOOTH/Xdffb3/M10_g N_VDD_XBOOTH/Xdffb3/M10_s
+ N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXBOOTH/Xsel23/M15 N_XBOOTH/XSEL23/N004_XBOOTH/Xsel23/M15_d
+ N_XBOOTH/XSEL23/B_XBOOTH/Xsel23/M15_g N_XBOOTH/XSEL23/N003_XBOOTH/Xsel23/M15_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel13/M15 N_XBOOTH/XSEL13/N004_XBOOTH/Xsel13/M15_d
+ N_XBOOTH/XSEL13/B_XBOOTH/Xsel13/M15_g N_XBOOTH/XSEL13/N003_XBOOTH/Xsel13/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel03/M15 N_XBOOTH/XSEL03/N004_XBOOTH/Xsel03/M15_d
+ N_XBOOTH/XSEL03/B_XBOOTH/Xsel03/M15_g N_XBOOTH/XSEL03/N003_XBOOTH/Xsel03/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mX02/xd29/M4 N_X02/XD29/N1_X02/xd29/M4_d N_CLK_X02/xd29/M4_g N_VDD_X02/xd29/M4_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa76/M5 N_XADDER/XA76/N002_XADDER/Xa76/M5_d N_XADDER/P6_XADDER/Xa76/M5_g
+ N_XADDER/XA76/N001_XADDER/Xa76/M5_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=4.444e-13 AS=6.16e-14 PD=2.46e-06 PS=2.8e-07
mXCSA/X_LV3_FA3/M3 N_XCSA/X_LV3_FA3/N001_XCSA/X_LV3_FA3/M3_d
+ N_XCSA/LV2_C[5]_XCSA/X_LV3_FA3/M3_g N_VDD_XCSA/X_LV3_FA3/M3_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA3/M1 N_XCSA/X_LV3_FA3/P001_XCSA/X_LV3_FA3/M1_d
+ N_XCSA/LV2_C[5]_XCSA/X_LV3_FA3/M1_g N_VDD_XCSA/X_LV3_FA3/M1_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA3/M10 N_XCSA/X_LV3_FA3/P002_XCSA/X_LV3_FA3/M10_d
+ N_XCSA/LV2_C[5]_XCSA/X_LV3_FA3/M10_g N_VDD_XCSA/X_LV3_FA3/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA3/M7 N_XCSA/X_LV3_FA3/N002_XCSA/X_LV3_FA3/M7_d
+ N_XCSA/LV2_C[5]_XCSA/X_LV3_FA3/M7_g N_VDD_XCSA/X_LV3_FA3/M7_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV1_FA3/M9 N_XCSA/X_LV1_FA3/_SUM_XCSA/X_LV1_FA3/M9_d
+ N_XCSA/X_LV1_FA3/_COUT_XCSA/X_LV1_FA3/M9_g
+ N_XCSA/X_LV1_FA3/N002_XCSA/X_LV1_FA3/M9_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXADDER/Xa66/Xao1/M12 N_XADDER/XA66/XAO1/N003_XADDER/Xa66/Xao1/M12_d
+ N_XADDER/P6_XADDER/Xa66/Xao1/M12_g N_VDD_XADDER/Xa66/Xao1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.288e-13 AS=1.474e-13
+ PD=1.48e-06 PS=6.7e-07
mXCSA/X_LV2_HA5/M13 N_XCSA/LV2_C[8]_XCSA/X_LV2_HA5/M13_d
+ N_XCSA/X_LV2_HA5/N001_XCSA/X_LV2_HA5/M13_g N_VDD_XCSA/X_LV2_HA5/M13_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA5/X_xor/M4 N_XCSA/LV2_S[7]_XCSA/X_LV2_HA5/X_xor/M4_d
+ N_XCSA/X_LV2_HA5/X_XOR/N002_XCSA/X_LV2_HA5/X_xor/M4_g
+ N_VDD_XCSA/X_LV2_HA5/X_xor/M4_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa76/M6 N_XADDER/XA76/N001_XADDER/Xa76/M6_d
+ N_XADDER/GX5[0]_XADDER/Xa76/M6_g N_VDD_XADDER/Xa76/M6_s N_VDD_XADDER/Xa72/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa5/M4 N_XCSA/XDFFA5/N1_XCSA/Xdffa5/M4_d N_CLK_XCSA/Xdffa5/M4_g
+ N_VDD_XCSA/Xdffa5/M4_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa18/M4 N_XCSA/XDFFA18/N1_XCSA/Xdffa18/M4_d N_CLK_XCSA/Xdffa18/M4_g
+ N_VDD_XCSA/Xdffa18/M4_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mX02/xd29/M7 N_X02/XD29/N3_X02/xd29/M7_d N_X02/XD29/N1_X02/xd29/M7_g
+ N_VDD_X02/xd29/M7_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA3/M28 N_XCSA/LV1_C[8]_XCSA/X_LV1_FA3/M28_d
+ N_XCSA/X_LV1_FA3/_COUT_XCSA/X_LV1_FA3/M28_g N_VDD_XCSA/X_LV1_FA3/M28_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa17/Xyb3/M36 N_XADDER/XA17/XYB3/N008_XADDER/Xa17/Xyb3/M36_d
+ N_XADDER/XA17/T1_XADDER/Xa17/Xyb3/M36_g
+ N_XADDER/XA17/XYB3/N007_XADDER/Xa17/Xyb3/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXADDER/Xa08/Xrb2/M4 N_XADDER/P7_XADDER/Xa08/Xrb2/M4_d
+ N_XADDER/XA08/XRB2/N002_XADDER/Xa08/Xrb2/M4_g N_VDD_XADDER/Xa08/Xrb2/M4_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel23/M14 N_PP2[3]_XBOOTH/Xsel23/M14_d
+ N_XBOOTH/XSEL23/N004_XBOOTH/Xsel23/M14_g N_VDD_XBOOTH/Xsel23/M14_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel13/M14 N_PP1[3]_XBOOTH/Xsel13/M14_d
+ N_XBOOTH/XSEL13/N004_XBOOTH/Xsel13/M14_g N_VDD_XBOOTH/Xsel13/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel03/M14 N_PP0[3]_XBOOTH/Xsel03/M14_d
+ N_XBOOTH/XSEL03/N004_XBOOTH/Xsel03/M14_g N_VDD_XBOOTH/Xsel03/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa5/M7 N_XCSA/XDFFA5/N3_XCSA/Xdffa5/M7_d
+ N_XCSA/XDFFA5/N1_XCSA/Xdffa5/M7_g N_VDD_XCSA/Xdffa5/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa18/M7 N_XCSA/XDFFA18/N3_XCSA/Xdffa18/M7_d
+ N_XCSA/XDFFA18/N1_XCSA/Xdffa18/M7_g N_VDD_XCSA/Xdffa18/M7_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa17/Xyb3/M35 N_XADDER/XA17/XYB3/N007_XADDER/Xa17/Xyb3/M35_d
+ N_XADDER/G7_XADDER/Xa17/Xyb3/M35_g N_VDD_XADDER/Xa17/Xyb3/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXCSA/X_LV1_FA3/M27 N_XCSA/LV1_S[7]_XCSA/X_LV1_FA3/M27_d
+ N_XCSA/X_LV1_FA3/_SUM_XCSA/X_LV1_FA3/M27_g N_VDD_XCSA/X_LV1_FA3/M27_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXCSA/X_LV3_FA4/M27 N_XCSA/LV3_S[6]_XCSA/X_LV3_FA4/M27_d
+ N_XCSA/X_LV3_FA4/_SUM_XCSA/X_LV3_FA4/M27_g N_VDD_XCSA/X_LV3_FA4/M27_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa66/Xao1/Xand1/M15 N_VDD_XADDER/Xa66/Xao1/Xand1/M15_d
+ N_XADDER/XA66/XAO1/N003_XADDER/Xa66/Xao1/Xand1/M15_g
+ N_XADDER/XA66/OUT1_XADDER/Xa66/Xao1/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd29/M10 N_OUT[8]_X02/xd29/M10_d N_X02/XD29/N3_X02/xd29/M10_g
+ N_VDD_X02/xd29/M10_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa17/Xyb3/Xor1/M15 N_VDD_XADDER/Xa17/Xyb3/Xor1/M15_d
+ N_XADDER/XA17/XYB3/N008_XADDER/Xa17/Xyb3/Xor1/M15_g
+ N_XADDER/GG7_XADDER/Xa17/Xyb3/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mXCSA/X_LV3_FA4/M28 N_XCSA/LV3_C[7]_XCSA/X_LV3_FA4/M28_d
+ N_XCSA/X_LV3_FA4/_COUT_XCSA/X_LV3_FA4/M28_g N_VDD_XCSA/X_LV3_FA4/M28_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa78/M4 N_OUT1[8]_XADDER/Xa78/M4_d N_XADDER/XA78/N002_XADDER/Xa78/M4_g
+ N_VDD_XADDER/Xa78/M4_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa08/Xrb2/M5 N_XADDER/XA08/XRB2/N001_XADDER/Xa08/Xrb2/M5_d
+ N_C[7]_XADDER/Xa08/Xrb2/M5_g N_VDD_XADDER/Xa08/Xrb2/M5_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.904e-13
+ PD=2.8e-07 PS=1.76e-06
mXCSA/Xdffa5/M10 N_C[6]_XCSA/Xdffa5/M10_d N_XCSA/XDFFA5/N3_XCSA/Xdffa5/M10_g
+ N_VDD_XCSA/Xdffa5/M10_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa18/M10 N_S[6]_XCSA/Xdffa18/M10_d N_XCSA/XDFFA18/N3_XCSA/Xdffa18/M10_g
+ N_VDD_XCSA/Xdffa18/M10_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA4/M9 N_XCSA/X_LV3_FA4/_SUM_XCSA/X_LV3_FA4/M9_d
+ N_XCSA/X_LV3_FA4/_COUT_XCSA/X_LV3_FA4/M9_g
+ N_XCSA/X_LV3_FA4/N002_XCSA/X_LV3_FA4/M9_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXADDER/Xa08/Xrb2/M6 N_XADDER/XA08/XRB2/N002_XADDER/Xa08/Xrb2/M6_d
+ N_S[7]_XADDER/Xa08/Xrb2/M6_g N_XADDER/XA08/XRB2/N001_XADDER/Xa08/Xrb2/M6_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa66/Xao2/M36 N_XADDER/XA66/XAO2/N008_XADDER/Xa66/Xao2/M36_d
+ N_XADDER/XA66/OUT1_XADDER/Xa66/Xao2/M36_g
+ N_XADDER/XA66/XAO2/N007_XADDER/Xa66/Xao2/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXBOOTH/Xsel24/M8 N_XBOOTH/XSEL24/N002_XBOOTH/Xsel24/M8_d
+ N_XBOOTH/B_D[3]_XBOOTH/Xsel24/M8_g N_noxref_1683_XBOOTH/Xsel24/M8_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel14/M8 N_XBOOTH/XSEL14/N002_XBOOTH/Xsel14/M8_d
+ N_XBOOTH/B_D[3]_XBOOTH/Xsel14/M8_g N_noxref_1684_XBOOTH/Xsel14/M8_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel04/M8 N_XBOOTH/XSEL04/N002_XBOOTH/Xsel04/M8_d
+ N_XBOOTH/B_D[3]_XBOOTH/Xsel04/M8_g N_noxref_1685_XBOOTH/Xsel04/M8_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mX02/xd210/M1 N_X02/XD210/P001_X02/xd210/M1_d N_OUT1[9]_X02/xd210/M1_g
+ N_VDD_X02/xd210/M1_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14
+ AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV1_FA4/M3 N_XCSA/X_LV1_FA4/N001_XCSA/X_LV1_FA4/M3_d
+ N_PP0[6]_XCSA/X_LV1_FA4/M3_g N_VDD_XCSA/X_LV1_FA4/M3_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV1_FA4/M1 N_XCSA/X_LV1_FA4/P001_XCSA/X_LV1_FA4/M1_d
+ N_PP0[6]_XCSA/X_LV1_FA4/M1_g N_VDD_XCSA/X_LV1_FA4/M1_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV1_FA4/M10 N_XCSA/X_LV1_FA4/P002_XCSA/X_LV1_FA4/M10_d
+ N_PP0[6]_XCSA/X_LV1_FA4/M10_g N_VDD_XCSA/X_LV1_FA4/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV1_FA4/M7 N_XCSA/X_LV1_FA4/N002_XCSA/X_LV1_FA4/M7_d
+ N_PP0[6]_XCSA/X_LV1_FA4/M7_g N_VDD_XCSA/X_LV1_FA4/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA4/M5 N_XCSA/X_LV3_FA4/_COUT_XCSA/X_LV3_FA4/M5_d
+ N_CACC[6]_XCSA/X_LV3_FA4/M5_g N_XCSA/X_LV3_FA4/N001_XCSA/X_LV3_FA4/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA4/M12 N_XCSA/X_LV3_FA4/_SUM_XCSA/X_LV3_FA4/M12_d
+ N_CACC[6]_XCSA/X_LV3_FA4/M12_g N_XCSA/X_LV3_FA4/P003_XCSA/X_LV3_FA4/M12_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA4/M6 N_XCSA/X_LV3_FA4/N002_XCSA/X_LV3_FA4/M6_d
+ N_CACC[6]_XCSA/X_LV3_FA4/M6_g N_VDD_XCSA/X_LV3_FA4/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV2_HA6/M9 N_XCSA/X_LV2_HA6/N001_XCSA/X_LV2_HA6/M9_d
+ N_XCSA/LV1_C[8]_XCSA/X_LV2_HA6/M9_g N_VDD_XCSA/X_LV2_HA6/M9_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA6/X_xor/M6 N_XCSA/X_LV2_HA6/X_XOR/N001_XCSA/X_LV2_HA6/X_xor/M6_d
+ N_XCSA/LV1_C[8]_XCSA/X_LV2_HA6/X_xor/M6_g N_VDD_XCSA/X_LV2_HA6/X_xor/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mX02/xd210/M2 N_X02/XD210/N0_X02/xd210/M2_d N_CLK_X02/xd210/M2_g
+ N_X02/XD210/P001_X02/xd210/M2_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa66/Xao2/M35 N_XADDER/XA66/XAO2/N007_XADDER/Xa66/Xao2/M35_d
+ N_XADDER/G6_XADDER/Xa66/Xao2/M35_g N_VDD_XADDER/Xa66/Xao2/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXBOOTH/Xsel24/M6 N_XBOOTH/XSEL24/N002_XBOOTH/Xsel24/M6_d
+ N_XBOOTH/D2_XBOOTH/Xsel24/M6_g N_noxref_1683_XBOOTH/Xsel24/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel14/M6 N_XBOOTH/XSEL14/N002_XBOOTH/Xsel14/M6_d
+ N_XBOOTH/D1_XBOOTH/Xsel14/M6_g N_noxref_1684_XBOOTH/Xsel14/M6_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel04/M6 N_XBOOTH/XSEL04/N002_XBOOTH/Xsel04/M6_d
+ N_XBOOTH/D0_XBOOTH/Xsel04/M6_g N_noxref_1685_XBOOTH/Xsel04/M6_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xdffb4/M1 N_XBOOTH/XDFFB4/P001_XBOOTH/Xdffb4/M1_d
+ N_B[4]_XBOOTH/Xdffb4/M1_g N_VDD_XBOOTH/Xdffb4/M1_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=7.7e-14 AS=2.695e-13 PD=2.8e-07 PS=1.53e-06
mXCSA/Xdffa6/M1 N_XCSA/XDFFA6/P001_XCSA/Xdffa6/M1_d
+ N_XCSA/LV3_C[7]_XCSA/Xdffa6/M1_g N_VDD_XCSA/Xdffa6/M1_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa19/M1 N_XCSA/XDFFA19/P001_XCSA/Xdffa19/M1_d
+ N_XCSA/LV3_S[7]_XCSA/Xdffa19/M1_g N_VDD_XCSA/Xdffa19/M1_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV1_FA4/M4 N_XCSA/X_LV1_FA4/N001_XCSA/X_LV1_FA4/M4_d
+ N_PP1[6]_XCSA/X_LV1_FA4/M4_g N_VDD_XCSA/X_LV1_FA4/M4_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA4/M2 N_XCSA/X_LV1_FA4/_COUT_XCSA/X_LV1_FA4/M2_d
+ N_PP1[6]_XCSA/X_LV1_FA4/M2_g N_XCSA/X_LV1_FA4/P001_XCSA/X_LV1_FA4/M2_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV1_FA4/M11 N_XCSA/X_LV1_FA4/P003_XCSA/X_LV1_FA4/M11_d
+ N_PP1[6]_XCSA/X_LV1_FA4/M11_g N_XCSA/X_LV1_FA4/P002_XCSA/X_LV1_FA4/M11_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA4/M8 N_XCSA/X_LV1_FA4/N002_XCSA/X_LV1_FA4/M8_d
+ N_PP1[6]_XCSA/X_LV1_FA4/M8_g N_VDD_XCSA/X_LV1_FA4/M8_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV2_HA6/X_xor/M5 N_XCSA/X_LV2_HA6/X_XOR/N002_XCSA/X_LV2_HA6/X_xor/M5_d
+ N_XCSA/LV1_S[8]_XCSA/X_LV2_HA6/X_xor/M5_g
+ N_XCSA/X_LV2_HA6/X_XOR/N001_XCSA/X_LV2_HA6/X_xor/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa78/M5 N_XADDER/XA78/N002_XADDER/Xa78/M5_d N_XADDER/P8_XADDER/Xa78/M5_g
+ N_XADDER/XA78/N001_XADDER/Xa78/M5_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=4.444e-13 AS=6.16e-14 PD=2.46e-06 PS=2.8e-07
mXBOOTH/Xdffb4/M2 N_XBOOTH/XDFFB4/N0_XBOOTH/Xdffb4/M2_d N_CLK_XBOOTH/Xdffb4/M2_g
+ N_XBOOTH/XDFFB4/P001_XBOOTH/Xdffb4/M2_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=7.7e-14 PD=1.53e-06 PS=2.8e-07
mXCSA/X_LV3_FA4/M4 N_XCSA/X_LV3_FA4/N001_XCSA/X_LV3_FA4/M4_d
+ N_XCSA/LV2_S[6]_XCSA/X_LV3_FA4/M4_g N_VDD_XCSA/X_LV3_FA4/M4_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA4/M2 N_XCSA/X_LV3_FA4/_COUT_XCSA/X_LV3_FA4/M2_d
+ N_XCSA/LV2_S[6]_XCSA/X_LV3_FA4/M2_g N_XCSA/X_LV3_FA4/P001_XCSA/X_LV3_FA4/M2_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA4/M11 N_XCSA/X_LV3_FA4/P003_XCSA/X_LV3_FA4/M11_d
+ N_XCSA/LV2_S[6]_XCSA/X_LV3_FA4/M11_g
+ N_XCSA/X_LV3_FA4/P002_XCSA/X_LV3_FA4/M11_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA4/M8 N_XCSA/X_LV3_FA4/N002_XCSA/X_LV3_FA4/M8_d
+ N_XCSA/LV2_S[6]_XCSA/X_LV3_FA4/M8_g N_VDD_XCSA/X_LV3_FA4/M8_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mXADDER/Xa08/Xrb1/M12 N_XADDER/XA08/XRB1/N003_XADDER/Xa08/Xrb1/M12_d
+ N_S[7]_XADDER/Xa08/Xrb1/M12_g N_VDD_XADDER/Xa08/Xrb1/M12_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa6/M2 N_XCSA/XDFFA6/N0_XCSA/Xdffa6/M2_d N_CLK_XCSA/Xdffa6/M2_g
+ N_XCSA/XDFFA6/P001_XCSA/Xdffa6/M2_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa19/M2 N_XCSA/XDFFA19/N0_XCSA/Xdffa19/M2_d N_CLK_XCSA/Xdffa19/M2_g
+ N_XCSA/XDFFA19/P001_XCSA/Xdffa19/M2_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV2_HA6/M10 N_XCSA/X_LV2_HA6/N001_XCSA/X_LV2_HA6/M10_d
+ N_XCSA/LV1_S[8]_XCSA/X_LV2_HA6/M10_g N_VDD_XCSA/X_LV2_HA6/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel24/M7 N_noxref_1683_XBOOTH/Xsel24/M7_d
+ N_XBOOTH/S2_XBOOTH/Xsel24/M7_g N_VDD_XBOOTH/Xsel24/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel14/M7 N_noxref_1684_XBOOTH/Xsel14/M7_d
+ N_XBOOTH/S1_XBOOTH/Xsel14/M7_g N_VDD_XBOOTH/Xsel14/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel04/M7 N_noxref_1685_XBOOTH/Xsel04/M7_d
+ N_XBOOTH/S0_XBOOTH/Xsel04/M7_g N_VDD_XBOOTH/Xsel04/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXADDER/Xa66/Xao2/Xor1/M15 N_VDD_XADDER/Xa66/Xao2/Xor1/M15_d
+ N_XADDER/XA66/XAO2/N008_XADDER/Xa66/Xao2/Xor1/M15_g
+ N_XADDER/GX6[2]_XADDER/Xa66/Xao2/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mXADDER/Xa77/M6 N_XADDER/XA77/N001_XADDER/Xa77/M6_d
+ N_XADDER/GX6[2]_XADDER/Xa77/M6_g N_VDD_XADDER/Xa77/M6_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXADDER/Xa78/M6 N_XADDER/XA78/N001_XADDER/Xa78/M6_d
+ N_XADDER/GOUT7_XADDER/Xa78/M6_g N_VDD_XADDER/Xa78/M6_s N_VDD_XADDER/Xa72/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV1_FA4/M5 N_XCSA/X_LV1_FA4/_COUT_XCSA/X_LV1_FA4/M5_d
+ N_PP2[4]_XCSA/X_LV1_FA4/M5_g N_XCSA/X_LV1_FA4/N001_XCSA/X_LV1_FA4/M5_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV1_FA4/M12 N_XCSA/X_LV1_FA4/_SUM_XCSA/X_LV1_FA4/M12_d
+ N_PP2[4]_XCSA/X_LV1_FA4/M12_g N_XCSA/X_LV1_FA4/P003_XCSA/X_LV1_FA4/M12_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV1_FA4/M6 N_XCSA/X_LV1_FA4/N002_XCSA/X_LV1_FA4/M6_d
+ N_PP2[4]_XCSA/X_LV1_FA4/M6_g N_VDD_XCSA/X_LV1_FA4/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA4/M3 N_XCSA/X_LV3_FA4/N001_XCSA/X_LV3_FA4/M3_d
+ N_XCSA/LV2_C[6]_XCSA/X_LV3_FA4/M3_g N_VDD_XCSA/X_LV3_FA4/M3_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA4/M1 N_XCSA/X_LV3_FA4/P001_XCSA/X_LV3_FA4/M1_d
+ N_XCSA/LV2_C[6]_XCSA/X_LV3_FA4/M1_g N_VDD_XCSA/X_LV3_FA4/M1_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA4/M10 N_XCSA/X_LV3_FA4/P002_XCSA/X_LV3_FA4/M10_d
+ N_XCSA/LV2_C[6]_XCSA/X_LV3_FA4/M10_g N_VDD_XCSA/X_LV3_FA4/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA4/M7 N_XCSA/X_LV3_FA4/N002_XCSA/X_LV3_FA4/M7_d
+ N_XCSA/LV2_C[6]_XCSA/X_LV3_FA4/M7_g N_VDD_XCSA/X_LV3_FA4/M7_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXADDER/Xa77/M5 N_XADDER/XA77/N002_XADDER/Xa77/M5_d N_XADDER/P7_XADDER/Xa77/M5_g
+ N_XADDER/XA77/N001_XADDER/Xa77/M5_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=4.444e-13 AS=6.16e-14 PD=2.46e-06 PS=2.8e-07
mXADDER/Xa08/Xrb1/M11 N_XADDER/XA08/XRB1/N003_XADDER/Xa08/Xrb1/M11_d
+ N_C[7]_XADDER/Xa08/Xrb1/M11_g N_VDD_XADDER/Xa08/Xrb1/M11_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd210/M4 N_X02/XD210/N1_X02/xd210/M4_d N_CLK_X02/xd210/M4_g
+ N_VDD_X02/xd210/M4_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel24/M9 N_noxref_1683_XBOOTH/Xsel24/M9_d
+ N_XBOOTH/B_D[4]_XBOOTH/Xsel24/M9_g N_VDD_XBOOTH/Xsel24/M9_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel14/M9 N_noxref_1684_XBOOTH/Xsel14/M9_d
+ N_XBOOTH/B_D[4]_XBOOTH/Xsel14/M9_g N_VDD_XBOOTH/Xsel14/M9_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel04/M9 N_noxref_1685_XBOOTH/Xsel04/M9_d
+ N_XBOOTH/B_D[4]_XBOOTH/Xsel04/M9_g N_VDD_XBOOTH/Xsel04/M9_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA4/M9 N_XCSA/X_LV1_FA4/_SUM_XCSA/X_LV1_FA4/M9_d
+ N_XCSA/X_LV1_FA4/_COUT_XCSA/X_LV1_FA4/M9_g
+ N_XCSA/X_LV1_FA4/N002_XCSA/X_LV1_FA4/M9_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXBOOTH/Xdffb4/M4 N_XBOOTH/XDFFB4/N1_XBOOTH/Xdffb4/M4_d N_CLK_XBOOTH/Xdffb4/M4_g
+ N_VDD_XBOOTH/Xdffb4/M4_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07
+ AD=2.695e-13 AS=1.485e-13 PD=1.53e-06 PS=5.4e-07
mXCSA/Xdffa6/M4 N_XCSA/XDFFA6/N1_XCSA/Xdffa6/M4_d N_CLK_XCSA/Xdffa6/M4_g
+ N_VDD_XCSA/Xdffa6/M4_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa19/M4 N_XCSA/XDFFA19/N1_XCSA/Xdffa19/M4_d N_CLK_XCSA/Xdffa19/M4_g
+ N_VDD_XCSA/Xdffa19/M4_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV2_HA6/M13 N_XCSA/LV2_C[9]_XCSA/X_LV2_HA6/M13_d
+ N_XCSA/X_LV2_HA6/N001_XCSA/X_LV2_HA6/M13_g N_VDD_XCSA/X_LV2_HA6/M13_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA6/X_xor/M4 N_XCSA/LV2_S[8]_XCSA/X_LV2_HA6/X_xor/M4_d
+ N_XCSA/X_LV2_HA6/X_XOR/N002_XCSA/X_LV2_HA6/X_xor/M4_g
+ N_VDD_XCSA/X_LV2_HA6/X_xor/M4_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd210/M7 N_X02/XD210/N3_X02/xd210/M7_d N_X02/XD210/N1_X02/xd210/M7_g
+ N_VDD_X02/xd210/M7_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel24/M10 N_XBOOTH/XSEL24/B_XBOOTH/Xsel24/M10_d
+ N_XBOOTH/XSEL24/N002_XBOOTH/Xsel24/M10_g N_VDD_XBOOTH/Xsel24/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel14/M10 N_XBOOTH/XSEL14/B_XBOOTH/Xsel14/M10_d
+ N_XBOOTH/XSEL14/N002_XBOOTH/Xsel14/M10_g N_VDD_XBOOTH/Xsel14/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel04/M10 N_XBOOTH/XSEL04/B_XBOOTH/Xsel04/M10_d
+ N_XBOOTH/XSEL04/N002_XBOOTH/Xsel04/M10_g N_VDD_XBOOTH/Xsel04/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA4/M28 N_XCSA/LV1_C[9]_XCSA/X_LV1_FA4/M28_d
+ N_XCSA/X_LV1_FA4/_COUT_XCSA/X_LV1_FA4/M28_g N_VDD_XCSA/X_LV1_FA4/M28_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXBOOTH/Xdffb4/M7 N_XBOOTH/XDFFB4/N3_XBOOTH/Xdffb4/M7_d
+ N_XBOOTH/XDFFB4/N1_XBOOTH/Xdffb4/M7_g N_VDD_XBOOTH/Xdffb4/M7_s
+ N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA5/M27 N_XCSA/LV3_S[7]_XCSA/X_LV3_FA5/M27_d
+ N_XCSA/X_LV3_FA5/_SUM_XCSA/X_LV3_FA5/M27_g N_VDD_XCSA/X_LV3_FA5/M27_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa08/Xrb1/Xand1/M15 N_VDD_XADDER/Xa08/Xrb1/Xand1/M15_d
+ N_XADDER/XA08/XRB1/N003_XADDER/Xa08/Xrb1/Xand1/M15_g
+ N_XADDER/G7_XADDER/Xa08/Xrb1/Xand1/M15_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa6/M7 N_XCSA/XDFFA6/N3_XCSA/Xdffa6/M7_d
+ N_XCSA/XDFFA6/N1_XCSA/Xdffa6/M7_g N_VDD_XCSA/Xdffa6/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa19/M7 N_XCSA/XDFFA19/N3_XCSA/Xdffa19/M7_d
+ N_XCSA/XDFFA19/N1_XCSA/Xdffa19/M7_g N_VDD_XCSA/Xdffa19/M7_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa77/M4 N_OUT1[7]_XADDER/Xa77/M4_d N_XADDER/XA77/N002_XADDER/Xa77/M4_g
+ N_VDD_XADDER/Xa77/M4_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA4/M27 N_XCSA/LV1_S[8]_XCSA/X_LV1_FA4/M27_d
+ N_XCSA/X_LV1_FA4/_SUM_XCSA/X_LV1_FA4/M27_g N_VDD_XCSA/X_LV1_FA4/M27_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa68/Xao1/M11 N_XADDER/XA68/XAO1/N003_XADDER/Xa68/Xao1/M11_d
+ N_XADDER/GOUT7_XADDER/Xa68/Xao1/M11_g N_VDD_XADDER/Xa68/Xao1/M11_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.474e-13
+ PD=1.42e-06 PS=6.7e-07
mXCSA/X_LV3_FA5/M28 N_XCSA/LV3_C[8]_XCSA/X_LV3_FA5/M28_d
+ N_XCSA/X_LV3_FA5/_COUT_XCSA/X_LV3_FA5/M28_g N_VDD_XCSA/X_LV3_FA5/M28_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mX02/xd210/M10 N_OUT[9]_X02/xd210/M10_d N_X02/XD210/N3_X02/xd210/M10_g
+ N_VDD_X02/xd210/M10_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa59/Xao1/M11 N_XADDER/XA59/XAO1/N003_XADDER/Xa59/Xao1/M11_d
+ N_XADDER/GOUT7_XADDER/Xa59/Xao1/M11_g N_VDD_XADDER/Xa59/Xao1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.474e-13
+ PD=1.42e-06 PS=6.7e-07
mXBOOTH/Xdffb4/M10 N_XBOOTH/B_D[4]_XBOOTH/Xdffb4/M10_d
+ N_XBOOTH/XDFFB4/N3_XBOOTH/Xdffb4/M10_g N_VDD_XBOOTH/Xdffb4/M10_s
+ N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXCSA/X_LV3_FA5/M9 N_XCSA/X_LV3_FA5/_SUM_XCSA/X_LV3_FA5/M9_d
+ N_XCSA/X_LV3_FA5/_COUT_XCSA/X_LV3_FA5/M9_g
+ N_XCSA/X_LV3_FA5/N002_XCSA/X_LV3_FA5/M9_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXBOOTH/Xsel24/M16 N_XBOOTH/XSEL24/N003_XBOOTH/Xsel24/M16_d
+ N_A_D[5]_XBOOTH/Xsel24/M16_g N_VDD_XBOOTH/Xsel24/M16_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel14/M16 N_XBOOTH/XSEL14/N003_XBOOTH/Xsel14/M16_d
+ N_A_D[3]_XBOOTH/Xsel14/M16_g N_VDD_XBOOTH/Xsel14/M16_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel04/M16 N_XBOOTH/XSEL04/N003_XBOOTH/Xsel04/M16_d
+ N_A_D[1]_XBOOTH/Xsel04/M16_g N_VDD_XBOOTH/Xsel04/M16_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXADDER/Xa68/Xao1/M12 N_XADDER/XA68/XAO1/N003_XADDER/Xa68/Xao1/M12_d
+ N_XADDER/P8_XADDER/Xa68/Xao1/M12_g N_VDD_XADDER/Xa68/Xao1/M12_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.288e-13 AS=1.474e-13
+ PD=1.48e-06 PS=6.7e-07
mXADDER/Xa09/Xrb2/M4 N_XADDER/P8_XADDER/Xa09/Xrb2/M4_d
+ N_XADDER/XA09/XRB2/N002_XADDER/Xa09/Xrb2/M4_g N_VDD_XADDER/Xa09/Xrb2/M4_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa6/M10 N_C[7]_XCSA/Xdffa6/M10_d N_XCSA/XDFFA6/N3_XCSA/Xdffa6/M10_g
+ N_VDD_XCSA/Xdffa6/M10_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa19/M10 N_S[7]_XCSA/Xdffa19/M10_d N_XCSA/XDFFA19/N3_XCSA/Xdffa19/M10_g
+ N_VDD_XCSA/Xdffa19/M10_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel24/M15 N_XBOOTH/XSEL24/N004_XBOOTH/Xsel24/M15_d
+ N_XBOOTH/XSEL24/B_XBOOTH/Xsel24/M15_g N_XBOOTH/XSEL24/N003_XBOOTH/Xsel24/M15_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel14/M15 N_XBOOTH/XSEL14/N004_XBOOTH/Xsel14/M15_d
+ N_XBOOTH/XSEL14/B_XBOOTH/Xsel14/M15_g N_XBOOTH/XSEL14/N003_XBOOTH/Xsel14/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel04/M15 N_XBOOTH/XSEL04/N004_XBOOTH/Xsel04/M15_d
+ N_XBOOTH/XSEL04/B_XBOOTH/Xsel04/M15_g N_XBOOTH/XSEL04/N003_XBOOTH/Xsel04/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa59/Xao1/M12 N_XADDER/XA59/XAO1/N003_XADDER/Xa59/Xao1/M12_d
+ N_XADDER/PP9_XADDER/Xa59/Xao1/M12_g N_VDD_XADDER/Xa59/Xao1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.288e-13 AS=1.474e-13
+ PD=1.48e-06 PS=6.7e-07
mXCSA/X_LV3_FA5/M5 N_XCSA/X_LV3_FA5/_COUT_XCSA/X_LV3_FA5/M5_d
+ N_CACC[7]_XCSA/X_LV3_FA5/M5_g N_XCSA/X_LV3_FA5/N001_XCSA/X_LV3_FA5/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA5/M12 N_XCSA/X_LV3_FA5/_SUM_XCSA/X_LV3_FA5/M12_d
+ N_CACC[7]_XCSA/X_LV3_FA5/M12_g N_XCSA/X_LV3_FA5/P003_XCSA/X_LV3_FA5/M12_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA5/M6 N_XCSA/X_LV3_FA5/N002_XCSA/X_LV3_FA5/M6_d
+ N_CACC[7]_XCSA/X_LV3_FA5/M6_g N_VDD_XCSA/X_LV3_FA5/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXADDER/Xa19/Xyb1/Xand1/M15 N_VDD_XADDER/Xa19/Xyb1/Xand1/M15_d
+ N_XADDER/XA19/XYB1/N003_XADDER/Xa19/Xyb1/Xand1/M15_g
+ N_XADDER/PP9_XADDER/Xa19/Xyb1/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd28/M1 N_X02/XD28/P001_X02/xd28/M1_d N_OUT1[7]_X02/xd28/M1_g
+ N_VDD_X02/xd28/M1_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14
+ AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV1_FA5/M3 N_XCSA/X_LV1_FA5/N001_XCSA/X_LV1_FA5/M3_d
+ N_XCSA/PP0_INVS_XCSA/X_LV1_FA5/M3_g N_VDD_XCSA/X_LV1_FA5/M3_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV1_FA5/M1 N_XCSA/X_LV1_FA5/P001_XCSA/X_LV1_FA5/M1_d
+ N_XCSA/PP0_INVS_XCSA/X_LV1_FA5/M1_g N_VDD_XCSA/X_LV1_FA5/M1_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV1_FA5/M10 N_XCSA/X_LV1_FA5/P002_XCSA/X_LV1_FA5/M10_d
+ N_XCSA/PP0_INVS_XCSA/X_LV1_FA5/M10_g N_VDD_XCSA/X_LV1_FA5/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV1_FA5/M7 N_XCSA/X_LV1_FA5/N002_XCSA/X_LV1_FA5/M7_d
+ N_XCSA/PP0_INVS_XCSA/X_LV1_FA5/M7_g N_VDD_XCSA/X_LV1_FA5/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mX02/xd28/M2 N_X02/XD28/N0_X02/xd28/M2_d N_CLK_X02/xd28/M2_g
+ N_X02/XD28/P001_X02/xd28/M2_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa68/Xao1/Xand1/M15 N_VDD_XADDER/Xa68/Xao1/Xand1/M15_d
+ N_XADDER/XA68/XAO1/N003_XADDER/Xa68/Xao1/Xand1/M15_g
+ N_XADDER/XA68/OUT1_XADDER/Xa68/Xao1/Xand1/M15_s N_VDD_XADDER/Xa72/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa7/M1 N_XCSA/XDFFA7/P001_XCSA/Xdffa7/M1_d
+ N_XCSA/LV3_C[8]_XCSA/Xdffa7/M1_g N_VDD_XCSA/Xdffa7/M1_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa20/M1 N_XCSA/XDFFA20/P001_XCSA/Xdffa20/M1_d
+ N_XCSA/LV3_S[8]_XCSA/Xdffa20/M1_g N_VDD_XCSA/Xdffa20/M1_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV3_FA5/M4 N_XCSA/X_LV3_FA5/N001_XCSA/X_LV3_FA5/M4_d
+ N_XCSA/LV2_S[7]_XCSA/X_LV3_FA5/M4_g N_VDD_XCSA/X_LV3_FA5/M4_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA5/M2 N_XCSA/X_LV3_FA5/_COUT_XCSA/X_LV3_FA5/M2_d
+ N_XCSA/LV2_S[7]_XCSA/X_LV3_FA5/M2_g N_XCSA/X_LV3_FA5/P001_XCSA/X_LV3_FA5/M2_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA5/M11 N_XCSA/X_LV3_FA5/P003_XCSA/X_LV3_FA5/M11_d
+ N_XCSA/LV2_S[7]_XCSA/X_LV3_FA5/M11_g
+ N_XCSA/X_LV3_FA5/P002_XCSA/X_LV3_FA5/M11_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA5/M8 N_XCSA/X_LV3_FA5/N002_XCSA/X_LV3_FA5/M8_d
+ N_XCSA/LV2_S[7]_XCSA/X_LV3_FA5/M8_g N_VDD_XCSA/X_LV3_FA5/M8_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mXBOOTH/Xsel24/M14 N_PP2[4]_XBOOTH/Xsel24/M14_d
+ N_XBOOTH/XSEL24/N004_XBOOTH/Xsel24/M14_g N_VDD_XBOOTH/Xsel24/M14_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel14/M14 N_PP1[4]_XBOOTH/Xsel14/M14_d
+ N_XBOOTH/XSEL14/N004_XBOOTH/Xsel14/M14_g N_VDD_XBOOTH/Xsel14/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel04/M14 N_PP0[4]_XBOOTH/Xsel04/M14_d
+ N_XBOOTH/XSEL04/N004_XBOOTH/Xsel04/M14_g N_VDD_XBOOTH/Xsel04/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa09/Xrb2/M5 N_XADDER/XA09/XRB2/N001_XADDER/Xa09/Xrb2/M5_d
+ N_C[8]_XADDER/Xa09/Xrb2/M5_g N_VDD_XADDER/Xa09/Xrb2/M5_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.904e-13
+ PD=2.8e-07 PS=1.76e-06
mXCSA/Xdffa7/M2 N_XCSA/XDFFA7/N0_XCSA/Xdffa7/M2_d N_CLK_XCSA/Xdffa7/M2_g
+ N_XCSA/XDFFA7/P001_XCSA/Xdffa7/M2_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa20/M2 N_XCSA/XDFFA20/N0_XCSA/Xdffa20/M2_d N_CLK_XCSA/Xdffa20/M2_g
+ N_XCSA/XDFFA20/P001_XCSA/Xdffa20/M2_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV1_FA5/M4 N_XCSA/X_LV1_FA5/N001_XCSA/X_LV1_FA5/M4_d
+ N_XCSA/PP1_INVS_XCSA/X_LV1_FA5/M4_g N_VDD_XCSA/X_LV1_FA5/M4_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA5/M2 N_XCSA/X_LV1_FA5/_COUT_XCSA/X_LV1_FA5/M2_d
+ N_XCSA/PP1_INVS_XCSA/X_LV1_FA5/M2_g N_XCSA/X_LV1_FA5/P001_XCSA/X_LV1_FA5/M2_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV1_FA5/M11 N_XCSA/X_LV1_FA5/P003_XCSA/X_LV1_FA5/M11_d
+ N_XCSA/PP1_INVS_XCSA/X_LV1_FA5/M11_g
+ N_XCSA/X_LV1_FA5/P002_XCSA/X_LV1_FA5/M11_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV1_FA5/M8 N_XCSA/X_LV1_FA5/N002_XCSA/X_LV1_FA5/M8_d
+ N_XCSA/PP1_INVS_XCSA/X_LV1_FA5/M8_g N_VDD_XCSA/X_LV1_FA5/M8_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV2_HA7/M9 N_XCSA/X_LV2_HA7/N001_XCSA/X_LV2_HA7/M9_d
+ N_XCSA/LV1_C[9]_XCSA/X_LV2_HA7/M9_g N_VDD_XCSA/X_LV2_HA7/M9_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA7/X_xor/M6 N_XCSA/X_LV2_HA7/X_XOR/N001_XCSA/X_LV2_HA7/X_xor/M6_d
+ N_XCSA/LV1_C[9]_XCSA/X_LV2_HA7/X_xor/M6_g N_VDD_XCSA/X_LV2_HA7/X_xor/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXADDER/Xa09/Xrb2/M6 N_XADDER/XA09/XRB2/N002_XADDER/Xa09/Xrb2/M6_d
+ N_S[8]_XADDER/Xa09/Xrb2/M6_g N_XADDER/XA09/XRB2/N001_XADDER/Xa09/Xrb2/M6_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa59/Xao1/Xand1/M15 N_VDD_XADDER/Xa59/Xao1/Xand1/M15_d
+ N_XADDER/XA59/XAO1/N003_XADDER/Xa59/Xao1/Xand1/M15_g
+ N_XADDER/XA59/OUT1_XADDER/Xa59/Xao1/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA5/M3 N_XCSA/X_LV3_FA5/N001_XCSA/X_LV3_FA5/M3_d
+ N_XCSA/LV2_C[7]_XCSA/X_LV3_FA5/M3_g N_VDD_XCSA/X_LV3_FA5/M3_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA5/M1 N_XCSA/X_LV3_FA5/P001_XCSA/X_LV3_FA5/M1_d
+ N_XCSA/LV2_C[7]_XCSA/X_LV3_FA5/M1_g N_VDD_XCSA/X_LV3_FA5/M1_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA5/M10 N_XCSA/X_LV3_FA5/P002_XCSA/X_LV3_FA5/M10_d
+ N_XCSA/LV2_C[7]_XCSA/X_LV3_FA5/M10_g N_VDD_XCSA/X_LV3_FA5/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA5/M7 N_XCSA/X_LV3_FA5/N002_XCSA/X_LV3_FA5/M7_d
+ N_XCSA/LV2_C[7]_XCSA/X_LV3_FA5/M7_g N_VDD_XCSA/X_LV3_FA5/M7_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXADDER/Xa19/Xyb1/M11 N_XADDER/XA19/XYB1/N003_XADDER/Xa19/Xyb1/M11_d
+ N_XADDER/P8_XADDER/Xa19/Xyb1/M11_g N_VDD_XADDER/Xa19/Xyb1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mXCSA/X_LV2_HA7/X_xor/M5 N_XCSA/X_LV2_HA7/X_XOR/N002_XCSA/X_LV2_HA7/X_xor/M5_d
+ N_XCSA/LV1_S[9]_XCSA/X_LV2_HA7/X_xor/M5_g
+ N_XCSA/X_LV2_HA7/X_XOR/N001_XCSA/X_LV2_HA7/X_xor/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV2_HA7/M10 N_XCSA/X_LV2_HA7/N001_XCSA/X_LV2_HA7/M10_d
+ N_XCSA/LV1_S[9]_XCSA/X_LV2_HA7/M10_g N_VDD_XCSA/X_LV2_HA7/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mX02/xd28/M4 N_X02/XD28/N1_X02/xd28/M4_d N_CLK_X02/xd28/M4_g N_VDD_X02/xd28/M4_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA5/M5 N_XCSA/X_LV1_FA5/_COUT_XCSA/X_LV1_FA5/M5_d
+ N_PP2[5]_XCSA/X_LV1_FA5/M5_g N_XCSA/X_LV1_FA5/N001_XCSA/X_LV1_FA5/M5_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV1_FA5/M12 N_XCSA/X_LV1_FA5/_SUM_XCSA/X_LV1_FA5/M12_d
+ N_PP2[5]_XCSA/X_LV1_FA5/M12_g N_XCSA/X_LV1_FA5/P003_XCSA/X_LV1_FA5/M12_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV1_FA5/M6 N_XCSA/X_LV1_FA5/N002_XCSA/X_LV1_FA5/M6_d
+ N_PP2[5]_XCSA/X_LV1_FA5/M6_g N_VDD_XCSA/X_LV1_FA5/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXADDER/Xa68/Xao2/M36 N_XADDER/XA68/XAO2/N008_XADDER/Xa68/Xao2/M36_d
+ N_XADDER/XA68/OUT1_XADDER/Xa68/Xao2/M36_g
+ N_XADDER/XA68/XAO2/N007_XADDER/Xa68/Xao2/M36_s N_VDD_XADDER/Xa72/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXADDER/Xa19/Xyb1/M12 N_XADDER/XA19/XYB1/N003_XADDER/Xa19/Xyb1/M12_d
+ N_XADDER/P9_XADDER/Xa19/Xyb1/M12_g N_VDD_XADDER/Xa19/Xyb1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa7/M4 N_XCSA/XDFFA7/N1_XCSA/Xdffa7/M4_d N_CLK_XCSA/Xdffa7/M4_g
+ N_VDD_XCSA/Xdffa7/M4_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa20/M4 N_XCSA/XDFFA20/N1_XCSA/Xdffa20/M4_d N_CLK_XCSA/Xdffa20/M4_g
+ N_VDD_XCSA/Xdffa20/M4_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mX02/xd28/M7 N_X02/XD28/N3_X02/xd28/M7_d N_X02/XD28/N1_X02/xd28/M7_g
+ N_VDD_X02/xd28/M7_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV1_FA5/M9 N_XCSA/X_LV1_FA5/_SUM_XCSA/X_LV1_FA5/M9_d
+ N_XCSA/X_LV1_FA5/_COUT_XCSA/X_LV1_FA5/M9_g
+ N_XCSA/X_LV1_FA5/N002_XCSA/X_LV1_FA5/M9_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXADDER/Xa68/Xao2/M35 N_XADDER/XA68/XAO2/N007_XADDER/Xa68/Xao2/M35_d
+ N_XADDER/G8_XADDER/Xa68/Xao2/M35_g N_VDD_XADDER/Xa68/Xao2/M35_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXADDER/Xa59/Xao2/M36 N_XADDER/XA59/XAO2/N008_XADDER/Xa59/Xao2/M36_d
+ N_XADDER/XA59/OUT1_XADDER/Xa59/Xao2/M36_g
+ N_XADDER/XA59/XAO2/N007_XADDER/Xa59/Xao2/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXCSA/X_LV3_FA6/M27 N_XCSA/LV3_S[8]_XCSA/X_LV3_FA6/M27_d
+ N_XCSA/X_LV3_FA6/_SUM_XCSA/X_LV3_FA6/M27_g N_VDD_XCSA/X_LV3_FA6/M27_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa09/Xrb1/M12 N_XADDER/XA09/XRB1/N003_XADDER/Xa09/Xrb1/M12_d
+ N_S[8]_XADDER/Xa09/Xrb1/M12_g N_VDD_XADDER/Xa09/Xrb1/M12_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel25/M8 N_XBOOTH/XSEL25/N002_XBOOTH/Xsel25/M8_d
+ N_XBOOTH/B_D[4]_XBOOTH/Xsel25/M8_g N_noxref_1727_XBOOTH/Xsel25/M8_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel15/M8 N_XBOOTH/XSEL15/N002_XBOOTH/Xsel15/M8_d
+ N_XBOOTH/B_D[4]_XBOOTH/Xsel15/M8_g N_noxref_1728_XBOOTH/Xsel15/M8_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel05/M8 N_XBOOTH/XSEL05/N002_XBOOTH/Xsel05/M8_d
+ N_XBOOTH/B_D[4]_XBOOTH/Xsel05/M8_g N_noxref_1729_XBOOTH/Xsel05/M8_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/Xdffa7/M7 N_XCSA/XDFFA7/N3_XCSA/Xdffa7/M7_d
+ N_XCSA/XDFFA7/N1_XCSA/Xdffa7/M7_g N_VDD_XCSA/Xdffa7/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa20/M7 N_XCSA/XDFFA20/N3_XCSA/Xdffa20/M7_d
+ N_XCSA/XDFFA20/N1_XCSA/Xdffa20/M7_g N_VDD_XCSA/Xdffa20/M7_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV2_HA7/M13 N_XCSA/LV2_C[10]_XCSA/X_LV2_HA7/M13_d
+ N_XCSA/X_LV2_HA7/N001_XCSA/X_LV2_HA7/M13_g N_VDD_XCSA/X_LV2_HA7/M13_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA7/X_xor/M4 N_XCSA/LV2_S[9]_XCSA/X_LV2_HA7/X_xor/M4_d
+ N_XCSA/X_LV2_HA7/X_XOR/N002_XCSA/X_LV2_HA7/X_xor/M4_g
+ N_VDD_XCSA/X_LV2_HA7/X_xor/M4_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA5/M28 N_XCSA/LV1_C[10]_XCSA/X_LV1_FA5/M28_d
+ N_XCSA/X_LV1_FA5/_COUT_XCSA/X_LV1_FA5/M28_g N_VDD_XCSA/X_LV1_FA5/M28_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXBOOTH/Xdffb5/M1 N_XBOOTH/XDFFB5/P001_XBOOTH/Xdffb5/M1_d
+ N_B[5]_XBOOTH/Xdffb5/M1_g N_VDD_XBOOTH/Xdffb5/M1_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=7.7e-14 AS=2.695e-13 PD=2.8e-07 PS=1.53e-06
mXADDER/Xa59/Xao2/M35 N_XADDER/XA59/XAO2/N007_XADDER/Xa59/Xao2/M35_d
+ N_XADDER/GG9_XADDER/Xa59/Xao2/M35_g N_VDD_XADDER/Xa59/Xao2/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXADDER/Xa68/Xao2/Xor1/M15 N_VDD_XADDER/Xa68/Xao2/Xor1/M15_d
+ N_XADDER/XA68/XAO2/N008_XADDER/Xa68/Xao2/Xor1/M15_g
+ N_XADDER/GX6[3]_XADDER/Xa68/Xao2/Xor1/M15_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mXADDER/Xa09/Xrb1/M11 N_XADDER/XA09/XRB1/N003_XADDER/Xa09/Xrb1/M11_d
+ N_C[8]_XADDER/Xa09/Xrb1/M11_g N_VDD_XADDER/Xa09/Xrb1/M11_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA6/M28 N_XCSA/LV3_C[9]_XCSA/X_LV3_FA6/M28_d
+ N_XCSA/X_LV3_FA6/_COUT_XCSA/X_LV3_FA6/M28_g N_VDD_XCSA/X_LV3_FA6/M28_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa19/Xyb2/M12 N_XADDER/XA19/XYB2/N003_XADDER/Xa19/Xyb2/M12_d
+ N_XADDER/P9_XADDER/Xa19/Xyb2/M12_g N_VDD_XADDER/Xa19/Xyb2/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel25/M6 N_XBOOTH/XSEL25/N002_XBOOTH/Xsel25/M6_d
+ N_XBOOTH/D2_XBOOTH/Xsel25/M6_g N_noxref_1727_XBOOTH/Xsel25/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel15/M6 N_XBOOTH/XSEL15/N002_XBOOTH/Xsel15/M6_d
+ N_XBOOTH/D1_XBOOTH/Xsel15/M6_g N_noxref_1728_XBOOTH/Xsel15/M6_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel05/M6 N_XBOOTH/XSEL05/N002_XBOOTH/Xsel05/M6_d
+ N_XBOOTH/D0_XBOOTH/Xsel05/M6_g N_noxref_1729_XBOOTH/Xsel05/M6_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xdffb5/M2 N_XBOOTH/XDFFB5/N0_XBOOTH/Xdffb5/M2_d N_CLK_XBOOTH/Xdffb5/M2_g
+ N_XBOOTH/XDFFB5/P001_XBOOTH/Xdffb5/M2_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07
+ W=5.5e-07 AD=2.695e-13 AS=7.7e-14 PD=1.53e-06 PS=2.8e-07
mX02/xd28/M10 N_OUT[7]_X02/xd28/M10_d N_X02/XD28/N3_X02/xd28/M10_g
+ N_VDD_X02/xd28/M10_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_FA5/M27 N_XCSA/LV1_S[9]_XCSA/X_LV1_FA5/M27_d
+ N_XCSA/X_LV1_FA5/_SUM_XCSA/X_LV1_FA5/M27_g N_VDD_XCSA/X_LV1_FA5/M27_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXCSA/X_LV3_FA6/M9 N_XCSA/X_LV3_FA6/_SUM_XCSA/X_LV3_FA6/M9_d
+ N_XCSA/X_LV3_FA6/_COUT_XCSA/X_LV3_FA6/M9_g
+ N_XCSA/X_LV3_FA6/N002_XCSA/X_LV3_FA6/M9_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXADDER/Xa59/Xao2/Xor1/M15 N_VDD_XADDER/Xa59/Xao2/Xor1/M15_d
+ N_XADDER/XA59/XAO2/N008_XADDER/Xa59/Xao2/Xor1/M15_g
+ N_XADDER/GX5[1]_XADDER/Xa59/Xao2/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mXADDER/Xa19/Xyb2/M11 N_XADDER/XA19/XYB2/N003_XADDER/Xa19/Xyb2/M11_d
+ N_XADDER/G8_XADDER/Xa19/Xyb2/M11_g N_VDD_XADDER/Xa19/Xyb2/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mXBOOTH/Xsel25/M7 N_noxref_1727_XBOOTH/Xsel25/M7_d
+ N_XBOOTH/S2_XBOOTH/Xsel25/M7_g N_VDD_XBOOTH/Xsel25/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel15/M7 N_noxref_1728_XBOOTH/Xsel15/M7_d
+ N_XBOOTH/S1_XBOOTH/Xsel15/M7_g N_VDD_XBOOTH/Xsel15/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel05/M7 N_noxref_1729_XBOOTH/Xsel05/M7_d
+ N_XBOOTH/S0_XBOOTH/Xsel05/M7_g N_VDD_XBOOTH/Xsel05/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXCSA/Xdffa7/M10 N_C[8]_XCSA/Xdffa7/M10_d N_XCSA/XDFFA7/N3_XCSA/Xdffa7/M10_g
+ N_VDD_XCSA/Xdffa7/M10_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa20/M10 N_S[8]_XCSA/Xdffa20/M10_d N_XCSA/XDFFA20/N3_XCSA/Xdffa20/M10_g
+ N_VDD_XCSA/Xdffa20/M10_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa09/Xrb1/Xand1/M15 N_VDD_XADDER/Xa09/Xrb1/Xand1/M15_d
+ N_XADDER/XA09/XRB1/N003_XADDER/Xa09/Xrb1/Xand1/M15_g
+ N_XADDER/G8_XADDER/Xa09/Xrb1/Xand1/M15_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA6/M5 N_XCSA/X_LV3_FA6/_COUT_XCSA/X_LV3_FA6/M5_d
+ N_CACC[8]_XCSA/X_LV3_FA6/M5_g N_XCSA/X_LV3_FA6/N001_XCSA/X_LV3_FA6/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA6/M12 N_XCSA/X_LV3_FA6/_SUM_XCSA/X_LV3_FA6/M12_d
+ N_CACC[8]_XCSA/X_LV3_FA6/M12_g N_XCSA/X_LV3_FA6/P003_XCSA/X_LV3_FA6/M12_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA6/M6 N_XCSA/X_LV3_FA6/N002_XCSA/X_LV3_FA6/M6_d
+ N_CACC[8]_XCSA/X_LV3_FA6/M6_g N_VDD_XCSA/X_LV3_FA6/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXBOOTH/Xsel25/M9 N_noxref_1727_XBOOTH/Xsel25/M9_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel25/M9_g N_VDD_XBOOTH/Xsel25/M9_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel15/M9 N_noxref_1728_XBOOTH/Xsel15/M9_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel15/M9_g N_VDD_XBOOTH/Xsel15/M9_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel05/M9 N_noxref_1729_XBOOTH/Xsel05/M9_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel05/M9_g N_VDD_XBOOTH/Xsel05/M9_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xdffb5/M4 N_XBOOTH/XDFFB5/N1_XBOOTH/Xdffb5/M4_d N_CLK_XBOOTH/Xdffb5/M4_g
+ N_VDD_XBOOTH/Xdffb5/M4_s N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07
+ AD=2.695e-13 AS=1.485e-13 PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA6/M4 N_XCSA/X_LV3_FA6/N001_XCSA/X_LV3_FA6/M4_d
+ N_XCSA/LV2_S[8]_XCSA/X_LV3_FA6/M4_g N_VDD_XCSA/X_LV3_FA6/M4_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA6/M2 N_XCSA/X_LV3_FA6/_COUT_XCSA/X_LV3_FA6/M2_d
+ N_XCSA/LV2_S[8]_XCSA/X_LV3_FA6/M2_g N_XCSA/X_LV3_FA6/P001_XCSA/X_LV3_FA6/M2_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA6/M11 N_XCSA/X_LV3_FA6/P003_XCSA/X_LV3_FA6/M11_d
+ N_XCSA/LV2_S[8]_XCSA/X_LV3_FA6/M11_g
+ N_XCSA/X_LV3_FA6/P002_XCSA/X_LV3_FA6/M11_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA6/M8 N_XCSA/X_LV3_FA6/N002_XCSA/X_LV3_FA6/M8_d
+ N_XCSA/LV2_S[8]_XCSA/X_LV3_FA6/M8_g N_VDD_XCSA/X_LV3_FA6/M8_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mXADDER/Xa19/Xyb2/Xand1/M15 N_VDD_XADDER/Xa19/Xyb2/Xand1/M15_d
+ N_XADDER/XA19/XYB2/N003_XADDER/Xa19/Xyb2/Xand1/M15_g
+ N_XADDER/XA19/T1_XADDER/Xa19/Xyb2/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xdffb5/M7 N_XBOOTH/XDFFB5/N3_XBOOTH/Xdffb5/M7_d
+ N_XBOOTH/XDFFB5/N1_XBOOTH/Xdffb5/M7_g N_VDD_XBOOTH/Xdffb5/M7_s
+ N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV2_HA8/M9 N_XCSA/X_LV2_HA8/N001_XCSA/X_LV2_HA8/M9_d
+ N_XCSA/LV1_C[10]_XCSA/X_LV2_HA8/M9_g N_VDD_XCSA/X_LV2_HA8/M9_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA8/X_xor/M6 N_XCSA/X_LV2_HA8/X_XOR/N001_XCSA/X_LV2_HA8/X_xor/M6_d
+ N_XCSA/LV1_C[10]_XCSA/X_LV2_HA8/X_xor/M6_g N_VDD_XCSA/X_LV2_HA8/X_xor/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV1_HA2/X_xor/M4 N_XCSA/LV1_S[10]_XCSA/X_LV1_HA2/X_xor/M4_d
+ N_XCSA/X_LV1_HA2/X_XOR/N002_XCSA/X_LV1_HA2/X_xor/M4_g
+ N_VDD_XCSA/X_LV1_HA2/X_xor/M4_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_HA2/M13 N_XCSA/LV1_C[11]_XCSA/X_LV1_HA2/M13_d
+ N_XCSA/X_LV1_HA2/N001_XCSA/X_LV1_HA2/M13_g N_VDD_XCSA/X_LV1_HA2/M13_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa79/M6 N_XADDER/XA79/N001_XADDER/Xa79/M6_d
+ N_XADDER/GX6[3]_XADDER/Xa79/M6_g N_VDD_XADDER/Xa79/M6_s N_VDD_XADDER/Xa72/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa8/M1 N_XCSA/XDFFA8/P001_XCSA/Xdffa8/M1_d
+ N_XCSA/LV3_C[9]_XCSA/Xdffa8/M1_g N_VDD_XCSA/Xdffa8/M1_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa21/M1 N_XCSA/XDFFA21/P001_XCSA/Xdffa21/M1_d
+ N_XCSA/LV3_S[9]_XCSA/Xdffa21/M1_g N_VDD_XCSA/Xdffa21/M1_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel25/M10 N_XBOOTH/XSEL25/B_XBOOTH/Xsel25/M10_d
+ N_XBOOTH/XSEL25/N002_XBOOTH/Xsel25/M10_g N_VDD_XBOOTH/Xsel25/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel15/M10 N_XBOOTH/XSEL15/B_XBOOTH/Xsel15/M10_d
+ N_XBOOTH/XSEL15/N002_XBOOTH/Xsel15/M10_g N_VDD_XBOOTH/Xsel15/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel05/M10 N_XBOOTH/XSEL05/B_XBOOTH/Xsel05/M10_d
+ N_XBOOTH/XSEL05/N002_XBOOTH/Xsel05/M10_g N_VDD_XBOOTH/Xsel05/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa010/Xrb2/M4 N_XADDER/P9_XADDER/Xa010/Xrb2/M4_d
+ N_XADDER/XA010/XRB2/N002_XADDER/Xa010/Xrb2/M4_g N_VDD_XADDER/Xa010/Xrb2/M4_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA8/X_xor/M5 N_XCSA/X_LV2_HA8/X_XOR/N002_XCSA/X_LV2_HA8/X_xor/M5_d
+ N_XCSA/LV1_S[10]_XCSA/X_LV2_HA8/X_xor/M5_g
+ N_XCSA/X_LV2_HA8/X_XOR/N001_XCSA/X_LV2_HA8/X_xor/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa79/M5 N_XADDER/XA79/N002_XADDER/Xa79/M5_d N_XADDER/P9_XADDER/Xa79/M5_g
+ N_XADDER/XA79/N001_XADDER/Xa79/M5_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=4.444e-13 AS=6.16e-14 PD=2.46e-06 PS=2.8e-07
mXCSA/X_LV3_FA6/M3 N_XCSA/X_LV3_FA6/N001_XCSA/X_LV3_FA6/M3_d
+ N_XCSA/LV2_C[8]_XCSA/X_LV3_FA6/M3_g N_VDD_XCSA/X_LV3_FA6/M3_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA6/M1 N_XCSA/X_LV3_FA6/P001_XCSA/X_LV3_FA6/M1_d
+ N_XCSA/LV2_C[8]_XCSA/X_LV3_FA6/M1_g N_VDD_XCSA/X_LV3_FA6/M1_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA6/M10 N_XCSA/X_LV3_FA6/P002_XCSA/X_LV3_FA6/M10_d
+ N_XCSA/LV2_C[8]_XCSA/X_LV3_FA6/M10_g N_VDD_XCSA/X_LV3_FA6/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA6/M7 N_XCSA/X_LV3_FA6/N002_XCSA/X_LV3_FA6/M7_d
+ N_XCSA/LV2_C[8]_XCSA/X_LV3_FA6/M7_g N_VDD_XCSA/X_LV3_FA6/M7_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/Xdffa8/M2 N_XCSA/XDFFA8/N0_XCSA/Xdffa8/M2_d N_CLK_XCSA/Xdffa8/M2_g
+ N_XCSA/XDFFA8/P001_XCSA/Xdffa8/M2_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa21/M2 N_XCSA/XDFFA21/N0_XCSA/Xdffa21/M2_d N_CLK_XCSA/Xdffa21/M2_g
+ N_XCSA/XDFFA21/P001_XCSA/Xdffa21/M2_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa211/Xyb1/Xand1/M15 N_VDD_XADDER/Xa211/Xyb1/Xand1/M15_d
+ N_XADDER/XA211/XYB1/N003_XADDER/Xa211/Xyb1/Xand1/M15_g
+ N_XADDER/PPP11_XADDER/Xa211/Xyb1/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA8/M10 N_XCSA/X_LV2_HA8/N001_XCSA/X_LV2_HA8/M10_d
+ N_XCSA/LV1_S[10]_XCSA/X_LV2_HA8/M10_g N_VDD_XCSA/X_LV2_HA8/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa19/Xyb3/M36 N_XADDER/XA19/XYB3/N008_XADDER/Xa19/Xyb3/M36_d
+ N_XADDER/XA19/T1_XADDER/Xa19/Xyb3/M36_g
+ N_XADDER/XA19/XYB3/N007_XADDER/Xa19/Xyb3/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXBOOTH/Xdffb5/M10 N_XBOOTH/B_D[5]_XBOOTH/Xdffb5/M10_d
+ N_XBOOTH/XDFFB5/N3_XBOOTH/Xdffb5/M10_g N_VDD_XBOOTH/Xdffb5/M10_s
+ N_VDD_XBOOTH/Xdffb0/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXCSA/X_LV1_HA2/M10 N_XCSA/X_LV1_HA2/N001_XCSA/X_LV1_HA2/M10_d
+ N_PP2[6]_XCSA/X_LV1_HA2/M10_g N_VDD_XCSA/X_LV1_HA2/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV1_HA2/X_xor/M5 N_XCSA/X_LV1_HA2/X_XOR/N002_XCSA/X_LV1_HA2/X_xor/M5_d
+ N_PP2[6]_XCSA/X_LV1_HA2/X_xor/M5_g
+ N_XCSA/X_LV1_HA2/X_XOR/N001_XCSA/X_LV1_HA2/X_xor/M5_s N_VDD_XBOOTH/Xdffa4/M1_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel25/M16 N_XBOOTH/XSEL25/N003_XBOOTH/Xsel25/M16_d
+ N_A_D[5]_XBOOTH/Xsel25/M16_g N_VDD_XBOOTH/Xsel25/M16_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel15/M16 N_XBOOTH/XSEL15/N003_XBOOTH/Xsel15/M16_d
+ N_A_D[3]_XBOOTH/Xsel15/M16_g N_VDD_XBOOTH/Xsel15/M16_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel05/M16 N_XBOOTH/XSEL05/N003_XBOOTH/Xsel05/M16_d
+ N_A_D[1]_XBOOTH/Xsel05/M16_g N_VDD_XBOOTH/Xsel05/M16_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa8/M4 N_XCSA/XDFFA8/N1_XCSA/Xdffa8/M4_d N_CLK_XCSA/Xdffa8/M4_g
+ N_VDD_XCSA/Xdffa8/M4_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA7/M27 N_XCSA/LV3_S[9]_XCSA/X_LV3_FA7/M27_d
+ N_XCSA/X_LV3_FA7/_SUM_XCSA/X_LV3_FA7/M27_g N_VDD_XCSA/X_LV3_FA7/M27_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXCSA/Xdffa21/M4 N_XCSA/XDFFA21/N1_XCSA/Xdffa21/M4_d N_CLK_XCSA/Xdffa21/M4_g
+ N_VDD_XCSA/Xdffa21/M4_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mX02/xd211/M1 N_X02/XD211/P001_X02/xd211/M1_d N_OUT1[10]_X02/xd211/M1_g
+ N_VDD_X02/xd211/M1_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14
+ AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXADDER/Xa19/Xyb3/M35 N_XADDER/XA19/XYB3/N007_XADDER/Xa19/Xyb3/M35_d
+ N_XADDER/G9_XADDER/Xa19/Xyb3/M35_g N_VDD_XADDER/Xa19/Xyb3/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXADDER/Xa010/Xrb2/M5 N_XADDER/XA010/XRB2/N001_XADDER/Xa010/Xrb2/M5_d
+ N_C[9]_XADDER/Xa010/Xrb2/M5_g N_VDD_XADDER/Xa010/Xrb2/M5_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.904e-13
+ PD=2.8e-07 PS=1.76e-06
mXCSA/X_LV2_HA8/M13 N_XCSA/LV2_C[11]_XCSA/X_LV2_HA8/M13_d
+ N_XCSA/X_LV2_HA8/N001_XCSA/X_LV2_HA8/M13_g N_VDD_XCSA/X_LV2_HA8/M13_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA8/X_xor/M4 N_XCSA/LV2_S[10]_XCSA/X_LV2_HA8/X_xor/M4_d
+ N_XCSA/X_LV2_HA8/X_XOR/N002_XCSA/X_LV2_HA8/X_xor/M4_g
+ N_VDD_XCSA/X_LV2_HA8/X_xor/M4_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV1_HA2/X_xor/M6 N_XCSA/X_LV1_HA2/X_XOR/N001_XCSA/X_LV1_HA2/X_xor/M6_d
+ N_VDD_XCSA/X_LV1_HA2/X_xor/M6_g N_VDD_XCSA/X_LV1_HA2/X_xor/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV1_HA2/M9 N_XCSA/X_LV1_HA2/N001_XCSA/X_LV1_HA2/M9_d
+ N_VDD_XCSA/X_LV1_HA2/M9_g N_VDD_XCSA/X_LV1_HA2/M9_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13 PD=5.4e-07 PS=1.44e-06
mXADDER/Xa211/Xyb1/M11 N_XADDER/XA211/XYB1/N003_XADDER/Xa211/Xyb1/M11_d
+ N_XADDER/PP9_XADDER/Xa211/Xyb1/M11_g N_VDD_XADDER/Xa211/Xyb1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mXBOOTH/Xsel25/M15 N_XBOOTH/XSEL25/N004_XBOOTH/Xsel25/M15_d
+ N_XBOOTH/XSEL25/B_XBOOTH/Xsel25/M15_g N_XBOOTH/XSEL25/N003_XBOOTH/Xsel25/M15_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel15/M15 N_XBOOTH/XSEL15/N004_XBOOTH/Xsel15/M15_d
+ N_XBOOTH/XSEL15/B_XBOOTH/Xsel15/M15_g N_XBOOTH/XSEL15/N003_XBOOTH/Xsel15/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel05/M15 N_XBOOTH/XSEL05/N004_XBOOTH/Xsel05/M15_d
+ N_XBOOTH/XSEL05/B_XBOOTH/Xsel05/M15_g N_XBOOTH/XSEL05/N003_XBOOTH/Xsel05/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa79/M4 N_OUT1[9]_XADDER/Xa79/M4_d N_XADDER/XA79/N002_XADDER/Xa79/M4_g
+ N_VDD_XADDER/Xa79/M4_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mX02/xd211/M2 N_X02/XD211/N0_X02/xd211/M2_d N_CLK_X02/xd211/M2_g
+ N_X02/XD211/P001_X02/xd211/M2_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa010/Xrb2/M6 N_XADDER/XA010/XRB2/N002_XADDER/Xa010/Xrb2/M6_d
+ N_S[9]_XADDER/Xa010/Xrb2/M6_g N_XADDER/XA010/XRB2/N001_XADDER/Xa010/Xrb2/M6_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa8/M7 N_XCSA/XDFFA8/N3_XCSA/Xdffa8/M7_d
+ N_XCSA/XDFFA8/N1_XCSA/Xdffa8/M7_g N_VDD_XCSA/Xdffa8/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa21/M7 N_XCSA/XDFFA21/N3_XCSA/Xdffa21/M7_d
+ N_XCSA/XDFFA21/N1_XCSA/Xdffa21/M7_g N_VDD_XCSA/Xdffa21/M7_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA7/M28 N_XCSA/LV3_C[10]_XCSA/X_LV3_FA7/M28_d
+ N_XCSA/X_LV3_FA7/_COUT_XCSA/X_LV3_FA7/M28_g N_VDD_XCSA/X_LV3_FA7/M28_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa19/Xyb3/Xor1/M15 N_VDD_XADDER/Xa19/Xyb3/Xor1/M15_d
+ N_XADDER/XA19/XYB3/N008_XADDER/Xa19/Xyb3/Xor1/M15_g
+ N_XADDER/GG9_XADDER/Xa19/Xyb3/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mXADDER/Xa211/Xyb1/M12 N_XADDER/XA211/XYB1/N003_XADDER/Xa211/Xyb1/M12_d
+ N_XADDER/PP11_XADDER/Xa211/Xyb1/M12_g N_VDD_XADDER/Xa211/Xyb1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA7/M9 N_XCSA/X_LV3_FA7/_SUM_XCSA/X_LV3_FA7/M9_d
+ N_XCSA/X_LV3_FA7/_COUT_XCSA/X_LV3_FA7/M9_g
+ N_XCSA/X_LV3_FA7/N002_XCSA/X_LV3_FA7/M9_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXBOOTH/Xsel25/M14 N_PP2[5]_XBOOTH/Xsel25/M14_d
+ N_XBOOTH/XSEL25/N004_XBOOTH/Xsel25/M14_g N_VDD_XBOOTH/Xsel25/M14_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel15/M14 N_PP1[5]_XBOOTH/Xsel15/M14_d
+ N_XBOOTH/XSEL15/N004_XBOOTH/Xsel15/M14_g N_VDD_XBOOTH/Xsel15/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel05/M14 N_PP0[5]_XBOOTH/Xsel05/M14_d
+ N_XBOOTH/XSEL05/N004_XBOOTH/Xsel05/M14_g N_VDD_XBOOTH/Xsel05/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mX02/xd211/M4 N_X02/XD211/N1_X02/xd211/M4_d N_CLK_X02/xd211/M4_g
+ N_VDD_X02/xd211/M4_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa8/M10 N_C[9]_XCSA/Xdffa8/M10_d N_XCSA/XDFFA8/N3_XCSA/Xdffa8/M10_g
+ N_VDD_XCSA/Xdffa8/M10_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa21/M10 N_S[9]_XCSA/Xdffa21/M10_d N_XCSA/XDFFA21/N3_XCSA/Xdffa21/M10_g
+ N_VDD_XCSA/Xdffa21/M10_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa411/Xao1/M11 N_XADDER/XA411/XAO1/N003_XADDER/Xa411/Xao1/M11_d
+ N_XADDER/GOUT7_XADDER/Xa411/Xao1/M11_g N_VDD_XADDER/Xa411/Xao1/M11_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.474e-13
+ PD=1.42e-06 PS=6.7e-07
mXCSA/X_LV3_FA7/M5 N_XCSA/X_LV3_FA7/_COUT_XCSA/X_LV3_FA7/M5_d
+ N_CACC[9]_XCSA/X_LV3_FA7/M5_g N_XCSA/X_LV3_FA7/N001_XCSA/X_LV3_FA7/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA7/M12 N_XCSA/X_LV3_FA7/_SUM_XCSA/X_LV3_FA7/M12_d
+ N_CACC[9]_XCSA/X_LV3_FA7/M12_g N_XCSA/X_LV3_FA7/P003_XCSA/X_LV3_FA7/M12_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA7/M6 N_XCSA/X_LV3_FA7/N002_XCSA/X_LV3_FA7/M6_d
+ N_CACC[9]_XCSA/X_LV3_FA7/M6_g N_VDD_XCSA/X_LV3_FA7/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXADDER/Xa010/Xrb1/M12 N_XADDER/XA010/XRB1/N003_XADDER/Xa010/Xrb1/M12_d
+ N_S[9]_XADDER/Xa010/Xrb1/M12_g N_VDD_XADDER/Xa010/Xrb1/M12_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa211/Xyb2/M12 N_XADDER/XA211/XYB2/N003_XADDER/Xa211/Xyb2/M12_d
+ N_XADDER/PP11_XADDER/Xa211/Xyb2/M12_g N_VDD_XADDER/Xa211/Xyb2/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd211/M7 N_X02/XD211/N3_X02/xd211/M7_d N_X02/XD211/N1_X02/xd211/M7_g
+ N_VDD_X02/xd211/M7_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXADDER/Xa010/Xrb1/M11 N_XADDER/XA010/XRB1/N003_XADDER/Xa010/Xrb1/M11_d
+ N_C[9]_XADDER/Xa010/Xrb1/M11_g N_VDD_XADDER/Xa010/Xrb1/M11_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA7/M4 N_XCSA/X_LV3_FA7/N001_XCSA/X_LV3_FA7/M4_d
+ N_XCSA/LV2_S[9]_XCSA/X_LV3_FA7/M4_g N_VDD_XCSA/X_LV3_FA7/M4_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA7/M2 N_XCSA/X_LV3_FA7/_COUT_XCSA/X_LV3_FA7/M2_d
+ N_XCSA/LV2_S[9]_XCSA/X_LV3_FA7/M2_g N_XCSA/X_LV3_FA7/P001_XCSA/X_LV3_FA7/M2_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA7/M11 N_XCSA/X_LV3_FA7/P003_XCSA/X_LV3_FA7/M11_d
+ N_XCSA/LV2_S[9]_XCSA/X_LV3_FA7/M11_g
+ N_XCSA/X_LV3_FA7/P002_XCSA/X_LV3_FA7/M11_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA7/M8 N_XCSA/X_LV3_FA7/N002_XCSA/X_LV3_FA7/M8_d
+ N_XCSA/LV2_S[9]_XCSA/X_LV3_FA7/M8_g N_VDD_XCSA/X_LV3_FA7/M8_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mXADDER/Xa411/Xao1/M12 N_XADDER/XA411/XAO1/N003_XADDER/Xa411/Xao1/M12_d
+ N_XADDER/PPP11_XADDER/Xa411/Xao1/M12_g N_VDD_XADDER/Xa411/Xao1/M12_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.288e-13 AS=1.474e-13
+ PD=1.48e-06 PS=6.7e-07
mXADDER/Xa610/Xao1/M11 N_XADDER/XA610/XAO1/N003_XADDER/Xa610/Xao1/M11_d
+ N_XADDER/GX5[1]_XADDER/Xa610/Xao1/M11_g N_VDD_XADDER/Xa610/Xao1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.474e-13
+ PD=1.42e-06 PS=6.7e-07
mXADDER/Xa211/Xyb2/M11 N_XADDER/XA211/XYB2/N003_XADDER/Xa211/Xyb2/M11_d
+ N_XADDER/GG9_XADDER/Xa211/Xyb2/M11_g N_VDD_XADDER/Xa211/Xyb2/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mXCSA/X_LV2_HA0/X_xor/M6 N_XCSA/X_LV2_HA0/X_XOR/N001_XCSA/X_LV2_HA0/X_xor/M6_d
+ N_PP0[0]_XCSA/X_LV2_HA0/X_xor/M6_g N_VDD_XCSA/X_LV2_HA0/X_xor/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV2_HA0/M9 N_XCSA/X_LV2_HA0/N001_XCSA/X_LV2_HA0/M9_d
+ N_PP0[0]_XCSA/X_LV2_HA0/M9_g N_VDD_XCSA/X_LV2_HA0/M9_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA9/M9 N_XCSA/X_LV2_HA9/N001_XCSA/X_LV2_HA9/M9_d
+ N_XCSA/LV1_C[11]_XCSA/X_LV2_HA9/M9_g N_VDD_XCSA/X_LV2_HA9/M9_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.2e-13
+ PD=5.4e-07 PS=1.44e-06
mXCSA/X_LV2_HA9/X_xor/M6 N_XCSA/X_LV2_HA9/X_XOR/N001_XCSA/X_LV2_HA9/X_xor/M6_d
+ N_XCSA/LV1_C[11]_XCSA/X_LV2_HA9/X_xor/M6_g N_VDD_XCSA/X_LV2_HA9/X_xor/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa9/M1 N_XCSA/XDFFA9/P001_XCSA/Xdffa9/M1_d
+ N_XCSA/LV3_C[10]_XCSA/Xdffa9/M1_g N_VDD_XCSA/Xdffa9/M1_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa22/M1 N_XCSA/XDFFA22/P001_XCSA/Xdffa22/M1_d
+ N_XCSA/LV3_S[10]_XCSA/Xdffa22/M1_g N_VDD_XCSA/Xdffa22/M1_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV3_FA7/M3 N_XCSA/X_LV3_FA7/N001_XCSA/X_LV3_FA7/M3_d
+ N_XCSA/LV2_C[9]_XCSA/X_LV3_FA7/M3_g N_VDD_XCSA/X_LV3_FA7/M3_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA7/M1 N_XCSA/X_LV3_FA7/P001_XCSA/X_LV3_FA7/M1_d
+ N_XCSA/LV2_C[9]_XCSA/X_LV3_FA7/M1_g N_VDD_XCSA/X_LV3_FA7/M1_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA7/M10 N_XCSA/X_LV3_FA7/P002_XCSA/X_LV3_FA7/M10_d
+ N_XCSA/LV2_C[9]_XCSA/X_LV3_FA7/M10_g N_VDD_XCSA/X_LV3_FA7/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA7/M7 N_XCSA/X_LV3_FA7/N002_XCSA/X_LV3_FA7/M7_d
+ N_XCSA/LV2_C[9]_XCSA/X_LV3_FA7/M7_g N_VDD_XCSA/X_LV3_FA7/M7_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXBOOTH/Xsel26/M8 N_XBOOTH/XSEL26/N002_XBOOTH/Xsel26/M8_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel26/M8_g N_XBOOTH/XSEL26/N001_XBOOTH/Xsel26/M8_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel16/M8 N_XBOOTH/XSEL16/N002_XBOOTH/Xsel16/M8_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel16/M8_g N_XBOOTH/XSEL16/N001_XBOOTH/Xsel16/M8_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXBOOTH/Xsel06/M8 N_XBOOTH/XSEL06/N002_XBOOTH/Xsel06/M8_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel06/M8_g N_XBOOTH/XSEL06/N001_XBOOTH/Xsel06/M8_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXCSA/X_LV2_HA0/X_xor/M5 N_XCSA/X_LV2_HA0/X_XOR/N002_XCSA/X_LV2_HA0/X_xor/M5_d
+ N_A_D[1]_XCSA/X_LV2_HA0/X_xor/M5_g
+ N_XCSA/X_LV2_HA0/X_XOR/N001_XCSA/X_LV2_HA0/X_xor/M5_s N_VDD_XBOOTH/Xdffa4/M1_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV2_HA9/X_xor/M5 N_XCSA/X_LV2_HA9/X_XOR/N002_XCSA/X_LV2_HA9/X_xor/M5_d
+ N_XCSA/PP2_INVS_XCSA/X_LV2_HA9/X_xor/M5_g
+ N_XCSA/X_LV2_HA9/X_XOR/N001_XCSA/X_LV2_HA9/X_xor/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXADDER/Xa610/Xao1/M12 N_XADDER/XA610/XAO1/N003_XADDER/Xa610/Xao1/M12_d
+ N_XADDER/P10_XADDER/Xa610/Xao1/M12_g N_VDD_XADDER/Xa610/Xao1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.288e-13 AS=1.474e-13
+ PD=1.48e-06 PS=6.7e-07
mXCSA/Xdffa9/M2 N_XCSA/XDFFA9/N0_XCSA/Xdffa9/M2_d N_CLK_XCSA/Xdffa9/M2_g
+ N_XCSA/XDFFA9/P001_XCSA/Xdffa9/M2_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa22/M2 N_XCSA/XDFFA22/N0_XCSA/Xdffa22/M2_d N_CLK_XCSA/Xdffa22/M2_g
+ N_XCSA/XDFFA22/P001_XCSA/Xdffa22/M2_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV2_HA0/M10 N_XCSA/X_LV2_HA0/N001_XCSA/X_LV2_HA0/M10_d
+ N_A_D[1]_XCSA/X_LV2_HA0/M10_g N_VDD_XCSA/X_LV2_HA0/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mX02/xd211/M10 N_OUT[10]_X02/xd211/M10_d N_X02/XD211/N3_X02/xd211/M10_g
+ N_VDD_X02/xd211/M10_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA9/M10 N_XCSA/X_LV2_HA9/N001_XCSA/X_LV2_HA9/M10_d
+ N_XCSA/PP2_INVS_XCSA/X_LV2_HA9/M10_g N_VDD_XCSA/X_LV2_HA9/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=2.156e-13
+ PD=5.4e-07 PS=1.42e-06
mXADDER/Xa010/Xrb1/Xand1/M15 N_VDD_XADDER/Xa010/Xrb1/Xand1/M15_d
+ N_XADDER/XA010/XRB1/N003_XADDER/Xa010/Xrb1/Xand1/M15_g
+ N_XADDER/G9_XADDER/Xa010/Xrb1/Xand1/M15_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa411/Xao1/Xand1/M15 N_VDD_XADDER/Xa411/Xao1/Xand1/M15_d
+ N_XADDER/XA411/XAO1/N003_XADDER/Xa411/Xao1/Xand1/M15_g
+ N_XADDER/XA411/OUT1_XADDER/Xa411/Xao1/Xand1/M15_s N_VDD_XADDER/Xa72/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel26/M6 N_XBOOTH/XSEL26/N002_XBOOTH/Xsel26/M6_d
+ N_XBOOTH/D2_XBOOTH/Xsel26/M6_g N_XBOOTH/XSEL26/N001_XBOOTH/Xsel26/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel16/M6 N_XBOOTH/XSEL16/N002_XBOOTH/Xsel16/M6_d
+ N_XBOOTH/D1_XBOOTH/Xsel16/M6_g N_XBOOTH/XSEL16/N001_XBOOTH/Xsel16/M6_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel06/M6 N_XBOOTH/XSEL06/N002_XBOOTH/Xsel06/M6_d
+ N_XBOOTH/D0_XBOOTH/Xsel06/M6_g N_XBOOTH/XSEL06/N001_XBOOTH/Xsel06/M6_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXADDER/Xa211/Xyb2/Xand1/M15 N_VDD_XADDER/Xa211/Xyb2/Xand1/M15_d
+ N_XADDER/XA211/XYB2/N003_XADDER/Xa211/Xyb2/Xand1/M15_g
+ N_XADDER/XA211/T1_XADDER/Xa211/Xyb2/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA8/M27 N_XCSA/LV3_S[10]_XCSA/X_LV3_FA8/M27_d
+ N_XCSA/X_LV3_FA8/_SUM_XCSA/X_LV3_FA8/M27_g N_VDD_XCSA/X_LV3_FA8/M27_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXBOOTH/Xsel26/M7 N_XBOOTH/XSEL26/N001_XBOOTH/Xsel26/M7_d
+ N_XBOOTH/S2_XBOOTH/Xsel26/M7_g N_VDD_XBOOTH/Xsel26/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel16/M7 N_XBOOTH/XSEL16/N001_XBOOTH/Xsel16/M7_d
+ N_XBOOTH/S1_XBOOTH/Xsel16/M7_g N_VDD_XBOOTH/Xsel16/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXBOOTH/Xsel06/M7 N_XBOOTH/XSEL06/N001_XBOOTH/Xsel06/M7_d
+ N_XBOOTH/S0_XBOOTH/Xsel06/M7_g N_VDD_XBOOTH/Xsel06/M7_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.188e-13 AS=1.188e-13
+ PD=5.4e-07 PS=5.4e-07
mXADDER/Xa610/Xao1/Xand1/M15 N_VDD_XADDER/Xa610/Xao1/Xand1/M15_d
+ N_XADDER/XA610/XAO1/N003_XADDER/Xa610/Xao1/Xand1/M15_g
+ N_XADDER/XA610/OUT1_XADDER/Xa610/Xao1/Xand1/M15_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa9/M4 N_XCSA/XDFFA9/N1_XCSA/Xdffa9/M4_d N_CLK_XCSA/Xdffa9/M4_g
+ N_VDD_XCSA/Xdffa9/M4_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa22/M4 N_XCSA/XDFFA22/N1_XCSA/Xdffa22/M4_d N_CLK_XCSA/Xdffa22/M4_g
+ N_VDD_XCSA/Xdffa22/M4_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV2_HA0/X_xor/M4 N_XCSA/LV2_S[0]_XCSA/X_LV2_HA0/X_xor/M4_d
+ N_XCSA/X_LV2_HA0/X_XOR/N002_XCSA/X_LV2_HA0/X_xor/M4_g
+ N_VDD_XCSA/X_LV2_HA0/X_xor/M4_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA0/M13 N_XCSA/LV2_C[1]_XCSA/X_LV2_HA0/M13_d
+ N_XCSA/X_LV2_HA0/N001_XCSA/X_LV2_HA0/M13_g N_VDD_XCSA/X_LV2_HA0/M13_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA9/M13 N_XCSA/LV2_C[12]_XCSA/X_LV2_HA9/M13_d
+ N_XCSA/X_LV2_HA9/N001_XCSA/X_LV2_HA9/M13_g N_VDD_XCSA/X_LV2_HA9/M13_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV2_HA9/X_xor/M4 N_XCSA/LV2_S[11]_XCSA/X_LV2_HA9/X_xor/M4_d
+ N_XCSA/X_LV2_HA9/X_XOR/N002_XCSA/X_LV2_HA9/X_xor/M4_g
+ N_VDD_XCSA/X_LV2_HA9/X_xor/M4_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa011/Xrb2/M4 N_XADDER/P10_XADDER/Xa011/Xrb2/M4_d
+ N_XADDER/XA011/XRB2/N002_XADDER/Xa011/Xrb2/M4_g N_VDD_XADDER/Xa011/Xrb2/M4_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa411/Xao2/M36 N_XADDER/XA411/XAO2/N008_XADDER/Xa411/Xao2/M36_d
+ N_XADDER/XA411/OUT1_XADDER/Xa411/Xao2/M36_g
+ N_XADDER/XA411/XAO2/N007_XADDER/Xa411/Xao2/M36_s N_VDD_XADDER/Xa72/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXBOOTH/Xsel26/M9 N_XBOOTH/XSEL26/N001_XBOOTH/Xsel26/M9_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel26/M9_g N_VDD_XBOOTH/Xsel26/M9_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel16/M9 N_XBOOTH/XSEL16/N001_XBOOTH/Xsel16/M9_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel16/M9_g N_VDD_XBOOTH/Xsel16/M9_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel06/M9 N_XBOOTH/XSEL06/N001_XBOOTH/Xsel06/M9_d
+ N_XBOOTH/B_D[5]_XBOOTH/Xsel06/M9_g N_VDD_XBOOTH/Xsel06/M9_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA8/M28 N_XCSA/LV3_C[11]_XCSA/X_LV3_FA8/M28_d
+ N_XCSA/X_LV3_FA8/_COUT_XCSA/X_LV3_FA8/M28_g N_VDD_XCSA/X_LV3_FA8/M28_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa211/Xyb3/M36 N_XADDER/XA211/XYB3/N008_XADDER/Xa211/Xyb3/M36_d
+ N_XADDER/XA211/T1_XADDER/Xa211/Xyb3/M36_g
+ N_XADDER/XA211/XYB3/N007_XADDER/Xa211/Xyb3/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXCSA/Xdffa9/M7 N_XCSA/XDFFA9/N3_XCSA/Xdffa9/M7_d
+ N_XCSA/XDFFA9/N1_XCSA/Xdffa9/M7_g N_VDD_XCSA/Xdffa9/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa22/M7 N_XCSA/XDFFA22/N3_XCSA/Xdffa22/M7_d
+ N_XCSA/XDFFA22/N1_XCSA/Xdffa22/M7_g N_VDD_XCSA/Xdffa22/M7_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA8/M9 N_XCSA/X_LV3_FA8/_SUM_XCSA/X_LV3_FA8/M9_d
+ N_XCSA/X_LV3_FA8/_COUT_XCSA/X_LV3_FA8/M9_g
+ N_XCSA/X_LV3_FA8/N002_XCSA/X_LV3_FA8/M9_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXADDER/Xa411/Xao2/M35 N_XADDER/XA411/XAO2/N007_XADDER/Xa411/Xao2/M35_d
+ N_XADDER/GGG11_XADDER/Xa411/Xao2/M35_g N_VDD_XADDER/Xa411/Xao2/M35_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXADDER/Xa610/Xao2/M36 N_XADDER/XA610/XAO2/N008_XADDER/Xa610/Xao2/M36_d
+ N_XADDER/XA610/OUT1_XADDER/Xa610/Xao2/M36_g
+ N_XADDER/XA610/XAO2/N007_XADDER/Xa610/Xao2/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mXADDER/Xa211/Xyb3/M35 N_XADDER/XA211/XYB3/N007_XADDER/Xa211/Xyb3/M35_d
+ N_XADDER/GG11_XADDER/Xa211/Xyb3/M35_g N_VDD_XADDER/Xa211/Xyb3/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXBOOTH/Xsel26/M10 N_XBOOTH/XSEL26/B_XBOOTH/Xsel26/M10_d
+ N_XBOOTH/XSEL26/N002_XBOOTH/Xsel26/M10_g N_VDD_XBOOTH/Xsel26/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel16/M10 N_XBOOTH/XSEL16/B_XBOOTH/Xsel16/M10_d
+ N_XBOOTH/XSEL16/N002_XBOOTH/Xsel16/M10_g N_VDD_XBOOTH/Xsel16/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel06/M10 N_XBOOTH/XSEL06/B_XBOOTH/Xsel06/M10_d
+ N_XBOOTH/XSEL06/N002_XBOOTH/Xsel06/M10_g N_VDD_XBOOTH/Xsel06/M10_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA8/M5 N_XCSA/X_LV3_FA8/_COUT_XCSA/X_LV3_FA8/M5_d
+ N_CACC[10]_XCSA/X_LV3_FA8/M5_g N_XCSA/X_LV3_FA8/N001_XCSA/X_LV3_FA8/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA8/M12 N_XCSA/X_LV3_FA8/_SUM_XCSA/X_LV3_FA8/M12_d
+ N_CACC[10]_XCSA/X_LV3_FA8/M12_g N_XCSA/X_LV3_FA8/P003_XCSA/X_LV3_FA8/M12_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA8/M6 N_XCSA/X_LV3_FA8/N002_XCSA/X_LV3_FA8/M6_d
+ N_CACC[10]_XCSA/X_LV3_FA8/M6_g N_VDD_XCSA/X_LV3_FA8/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXADDER/Xa411/Xao2/Xor1/M15 N_VDD_XADDER/Xa411/Xao2/Xor1/M15_d
+ N_XADDER/XA411/XAO2/N008_XADDER/Xa411/Xao2/Xor1/M15_g
+ N_XADDER/FG11_XADDER/Xa411/Xao2/Xor1/M15_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mXCSA/X_LV3_FA10/M3 N_XCSA/X_LV3_FA10/N001_XCSA/X_LV3_FA10/M3_d
+ N_XCSA/LV2_C[12]_XCSA/X_LV3_FA10/M3_g N_VDD_XCSA/X_LV3_FA10/M3_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA10/M1 N_XCSA/X_LV3_FA10/P001_XCSA/X_LV3_FA10/M1_d
+ N_XCSA/LV2_C[12]_XCSA/X_LV3_FA10/M1_g N_VDD_XCSA/X_LV3_FA10/M1_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA10/M10 N_XCSA/X_LV3_FA10/P002_XCSA/X_LV3_FA10/M10_d
+ N_XCSA/LV2_C[12]_XCSA/X_LV3_FA10/M10_g N_VDD_XCSA/X_LV3_FA10/M10_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA10/M7 N_XCSA/X_LV3_FA10/N002_XCSA/X_LV3_FA10/M7_d
+ N_XCSA/LV2_C[12]_XCSA/X_LV3_FA10/M7_g N_VDD_XCSA/X_LV3_FA10/M7_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXADDER/Xa011/Xrb2/M5 N_XADDER/XA011/XRB2/N001_XADDER/Xa011/Xrb2/M5_d
+ N_C[10]_XADDER/Xa011/Xrb2/M5_g N_VDD_XADDER/Xa011/Xrb2/M5_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.904e-13
+ PD=2.8e-07 PS=1.76e-06
mXADDER/Xa610/Xao2/M35 N_XADDER/XA610/XAO2/N007_XADDER/Xa610/Xao2/M35_d
+ N_XADDER/G10_XADDER/Xa610/Xao2/M35_g N_VDD_XADDER/Xa610/Xao2/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXCSA/Xdffa9/M10 N_C[10]_XCSA/Xdffa9/M10_d N_XCSA/XDFFA9/N3_XCSA/Xdffa9/M10_g
+ N_VDD_XCSA/Xdffa9/M10_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa22/M10 N_S[10]_XCSA/Xdffa22/M10_d
+ N_XCSA/XDFFA22/N3_XCSA/Xdffa22/M10_g N_VDD_XCSA/Xdffa22/M10_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa211/Xyb3/Xor1/M15 N_VDD_XADDER/Xa211/Xyb3/Xor1/M15_d
+ N_XADDER/XA211/XYB3/N008_XADDER/Xa211/Xyb3/Xor1/M15_g
+ N_XADDER/GGG11_XADDER/Xa211/Xyb3/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mXCSA/X_LV3_FA9/M7 N_XCSA/X_LV3_FA9/N002_XCSA/X_LV3_FA9/M7_d
+ N_XCSA/LV2_C[11]_XCSA/X_LV3_FA9/M7_g N_VDD_XCSA/X_LV3_FA9/M7_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA9/M10 N_XCSA/X_LV3_FA9/P002_XCSA/X_LV3_FA9/M10_d
+ N_XCSA/LV2_C[11]_XCSA/X_LV3_FA9/M10_g N_VDD_XCSA/X_LV3_FA9/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA9/M1 N_XCSA/X_LV3_FA9/P001_XCSA/X_LV3_FA9/M1_d
+ N_XCSA/LV2_C[11]_XCSA/X_LV3_FA9/M1_g N_VDD_XCSA/X_LV3_FA9/M1_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA9/M3 N_XCSA/X_LV3_FA9/N001_XCSA/X_LV3_FA9/M3_d
+ N_XCSA/LV2_C[11]_XCSA/X_LV3_FA9/M3_g N_VDD_XCSA/X_LV3_FA9/M3_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXADDER/Xa011/Xrb2/M6 N_XADDER/XA011/XRB2/N002_XADDER/Xa011/Xrb2/M6_d
+ N_S[10]_XADDER/Xa011/Xrb2/M6_g N_XADDER/XA011/XRB2/N001_XADDER/Xa011/Xrb2/M6_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV3_FA8/M4 N_XCSA/X_LV3_FA8/N001_XCSA/X_LV3_FA8/M4_d
+ N_XCSA/LV2_S[10]_XCSA/X_LV3_FA8/M4_g N_VDD_XCSA/X_LV3_FA8/M4_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA8/M2 N_XCSA/X_LV3_FA8/_COUT_XCSA/X_LV3_FA8/M2_d
+ N_XCSA/LV2_S[10]_XCSA/X_LV3_FA8/M2_g N_XCSA/X_LV3_FA8/P001_XCSA/X_LV3_FA8/M2_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA8/M11 N_XCSA/X_LV3_FA8/P003_XCSA/X_LV3_FA8/M11_d
+ N_XCSA/LV2_S[10]_XCSA/X_LV3_FA8/M11_g
+ N_XCSA/X_LV3_FA8/P002_XCSA/X_LV3_FA8/M11_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA8/M8 N_XCSA/X_LV3_FA8/N002_XCSA/X_LV3_FA8/M8_d
+ N_XCSA/LV2_S[10]_XCSA/X_LV3_FA8/M8_g N_VDD_XCSA/X_LV3_FA8/M8_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA10/M4 N_XCSA/X_LV3_FA10/N001_XCSA/X_LV3_FA10/M4_d
+ N_VDD_XCSA/X_LV3_FA10/M4_g N_VDD_XCSA/X_LV3_FA10/M4_s N_VDD_XBOOTH/Xdffa4/M1_b
+ P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA10/M2 N_XCSA/X_LV3_FA10/_COUT_XCSA/X_LV3_FA10/M2_d
+ N_VDD_XCSA/X_LV3_FA10/M2_g N_XCSA/X_LV3_FA10/P001_XCSA/X_LV3_FA10/M2_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA10/M11 N_XCSA/X_LV3_FA10/P003_XCSA/X_LV3_FA10/M11_d
+ N_VDD_XCSA/X_LV3_FA10/M11_g N_XCSA/X_LV3_FA10/P002_XCSA/X_LV3_FA10/M11_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA10/M8 N_XCSA/X_LV3_FA10/N002_XCSA/X_LV3_FA10/M8_d
+ N_VDD_XCSA/X_LV3_FA10/M8_g N_VDD_XCSA/X_LV3_FA10/M8_s N_VDD_XBOOTH/Xdffa4/M1_b
+ P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13 PD=5.4e-07 PS=5.9e-07
mXADDER/Xa610/Xao2/Xor1/M15 N_VDD_XADDER/Xa610/Xao2/Xor1/M15_d
+ N_XADDER/XA610/XAO2/N008_XADDER/Xa610/Xao2/Xor1/M15_g
+ N_XADDER/GX6[4]_XADDER/Xa610/Xao2/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
mXCSA/X_LV3_FA9/M8 N_XCSA/X_LV3_FA9/N002_XCSA/X_LV3_FA9/M8_d
+ N_XCSA/LV2_S[11]_XCSA/X_LV3_FA9/M8_g N_VDD_XCSA/X_LV3_FA9/M8_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=1.6225e-13
+ PD=5.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA9/M11 N_XCSA/X_LV3_FA9/P003_XCSA/X_LV3_FA9/M11_d
+ N_XCSA/LV2_S[11]_XCSA/X_LV3_FA9/M11_g
+ N_XCSA/X_LV3_FA9/P002_XCSA/X_LV3_FA9/M11_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13 PD=5.9e-07 PS=5.4e-07
mXCSA/X_LV3_FA9/M2 N_XCSA/X_LV3_FA9/_COUT_XCSA/X_LV3_FA9/M2_d
+ N_XCSA/LV2_S[11]_XCSA/X_LV3_FA9/M2_g N_XCSA/X_LV3_FA9/P001_XCSA/X_LV3_FA9/M2_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA9/M4 N_XCSA/X_LV3_FA9/N001_XCSA/X_LV3_FA9/M4_d
+ N_XCSA/LV2_S[11]_XCSA/X_LV3_FA9/M4_g N_VDD_XCSA/X_LV3_FA9/M4_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.6225e-13 AS=1.485e-13
+ PD=5.9e-07 PS=5.4e-07
mXBOOTH/Xsel26/M16 N_XBOOTH/XSEL26/N003_XBOOTH/Xsel26/M16_d
+ N_A_D[5]_XBOOTH/Xsel26/M16_g N_VDD_XBOOTH/Xsel26/M16_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel16/M16 N_XBOOTH/XSEL16/N003_XBOOTH/Xsel16/M16_d
+ N_A_D[3]_XBOOTH/Xsel16/M16_g N_VDD_XBOOTH/Xsel16/M16_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel06/M16 N_XBOOTH/XSEL06/N003_XBOOTH/Xsel06/M16_d
+ N_A_D[1]_XBOOTH/Xsel06/M16_g N_VDD_XBOOTH/Xsel06/M16_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mX02/xd212/M1 N_X02/XD212/P001_X02/xd212/M1_d N_OUT1[11]_X02/xd212/M1_g
+ N_VDD_X02/xd212/M1_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14
+ AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV3_FA8/M3 N_XCSA/X_LV3_FA8/N001_XCSA/X_LV3_FA8/M3_d
+ N_XCSA/LV2_C[10]_XCSA/X_LV3_FA8/M3_g N_VDD_XCSA/X_LV3_FA8/M3_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.485e-13
+ PD=1.53e-06 PS=5.4e-07
mXCSA/X_LV3_FA8/M1 N_XCSA/X_LV3_FA8/P001_XCSA/X_LV3_FA8/M1_d
+ N_XCSA/LV2_C[10]_XCSA/X_LV3_FA8/M1_g N_VDD_XCSA/X_LV3_FA8/M1_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA8/M10 N_XCSA/X_LV3_FA8/P002_XCSA/X_LV3_FA8/M10_d
+ N_XCSA/LV2_C[10]_XCSA/X_LV3_FA8/M10_g N_VDD_XCSA/X_LV3_FA8/M10_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA8/M7 N_XCSA/X_LV3_FA8/N002_XCSA/X_LV3_FA8/M7_d
+ N_XCSA/LV2_C[10]_XCSA/X_LV3_FA8/M7_g N_VDD_XCSA/X_LV3_FA8/M7_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.485e-13 AS=2.695e-13
+ PD=5.4e-07 PS=1.53e-06
mXCSA/X_LV3_FA10/M5 N_XCSA/X_LV3_FA10/_COUT_XCSA/X_LV3_FA10/M5_d
+ N_CACC[11]_XCSA/X_LV3_FA10/M5_g N_XCSA/X_LV3_FA10/N001_XCSA/X_LV3_FA10/M5_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA10/M12 N_XCSA/X_LV3_FA10/_SUM_XCSA/X_LV3_FA10/M12_d
+ N_CACC[11]_XCSA/X_LV3_FA10/M12_g N_XCSA/X_LV3_FA10/P003_XCSA/X_LV3_FA10/M12_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA10/M6 N_XCSA/X_LV3_FA10/N002_XCSA/X_LV3_FA10/M6_d
+ N_CACC[11]_XCSA/X_LV3_FA10/M6_g N_VDD_XCSA/X_LV3_FA10/M6_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/Xdffa10/M1 N_XCSA/XDFFA10/P001_XCSA/Xdffa10/M1_d
+ N_XCSA/LV3_C[11]_XCSA/Xdffa10/M1_g N_VDD_XCSA/Xdffa10/M1_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa23/M1 N_XCSA/XDFFA23/P001_XCSA/Xdffa23/M1_d
+ N_XCSA/LV3_S[11]_XCSA/Xdffa23/M1_g N_VDD_XCSA/Xdffa23/M1_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXBOOTH/Xsel26/M15 N_XBOOTH/XSEL26/N004_XBOOTH/Xsel26/M15_d
+ N_XBOOTH/XSEL26/B_XBOOTH/Xsel26/M15_g N_XBOOTH/XSEL26/N003_XBOOTH/Xsel26/M15_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel16/M15 N_XBOOTH/XSEL16/N004_XBOOTH/Xsel16/M15_d
+ N_XBOOTH/XSEL16/B_XBOOTH/Xsel16/M15_g N_XBOOTH/XSEL16/N003_XBOOTH/Xsel16/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mXBOOTH/Xsel06/M15 N_XBOOTH/XSEL06/N004_XBOOTH/Xsel06/M15_d
+ N_XBOOTH/XSEL06/B_XBOOTH/Xsel06/M15_g N_XBOOTH/XSEL06/N003_XBOOTH/Xsel06/M15_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mX02/xd212/M2 N_X02/XD212/N0_X02/xd212/M2_d N_CLK_X02/xd212/M2_g
+ N_X02/XD212/P001_X02/xd212/M2_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/X_LV3_FA9/M6 N_XCSA/X_LV3_FA9/N002_XCSA/X_LV3_FA9/M6_d
+ N_CACC[11]_XCSA/X_LV3_FA9/M6_g N_VDD_XCSA/X_LV3_FA9/M6_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=1.76e-13 AS=1.6225e-13
+ PD=6.4e-07 PS=5.9e-07
mXCSA/X_LV3_FA9/M12 N_XCSA/X_LV3_FA9/_SUM_XCSA/X_LV3_FA9/M12_d
+ N_CACC[11]_XCSA/X_LV3_FA9/M12_g N_XCSA/X_LV3_FA9/P003_XCSA/X_LV3_FA9/M12_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/X_LV3_FA9/M5 N_XCSA/X_LV3_FA9/_COUT_XCSA/X_LV3_FA9/M5_d
+ N_CACC[11]_XCSA/X_LV3_FA9/M5_g N_XCSA/X_LV3_FA9/N001_XCSA/X_LV3_FA9/M5_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.6225e-13
+ PD=1.53e-06 PS=5.9e-07
mXCSA/Xdffa10/M2 N_XCSA/XDFFA10/N0_XCSA/Xdffa10/M2_d N_CLK_XCSA/Xdffa10/M2_g
+ N_XCSA/XDFFA10/P001_XCSA/Xdffa10/M2_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa23/M2 N_XCSA/XDFFA23/N0_XCSA/Xdffa23/M2_d N_CLK_XCSA/Xdffa23/M2_g
+ N_XCSA/XDFFA23/P001_XCSA/Xdffa23/M2_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa011/Xrb1/M12 N_XADDER/XA011/XRB1/N003_XADDER/Xa011/Xrb1/M12_d
+ N_S[10]_XADDER/Xa011/Xrb1/M12_g N_VDD_XADDER/Xa011/Xrb1/M12_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA10/M9 N_XCSA/X_LV3_FA10/_SUM_XCSA/X_LV3_FA10/M9_d
+ N_XCSA/X_LV3_FA10/_COUT_XCSA/X_LV3_FA10/M9_g
+ N_XCSA/X_LV3_FA10/N002_XCSA/X_LV3_FA10/M9_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXADDER/Xa712/M6 N_XADDER/XA712/N001_XADDER/Xa712/M6_d
+ N_XADDER/FG11_XADDER/Xa712/M6_g N_VDD_XADDER/Xa712/M6_s N_VDD_XADDER/Xa72/M4_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXCSA/X_LV3_FA9/M9 N_XCSA/X_LV3_FA9/_SUM_XCSA/X_LV3_FA9/M9_d
+ N_XCSA/X_LV3_FA9/_COUT_XCSA/X_LV3_FA9/M9_g
+ N_XCSA/X_LV3_FA9/N002_XCSA/X_LV3_FA9/M9_s N_VDD_XACCXOR/X_xor2/M4_b P_18_G2
+ L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=1.76e-13 PD=1.53e-06 PS=6.4e-07
mXADDER/Xa111/Xyb1/Xand1/M15 N_VDD_XADDER/Xa111/Xyb1/Xand1/M15_d
+ N_XADDER/XA111/XYB1/N003_XADDER/Xa111/Xyb1/Xand1/M15_g
+ N_XADDER/PP11_XADDER/Xa111/Xyb1/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa011/Xrb1/M11 N_XADDER/XA011/XRB1/N003_XADDER/Xa011/Xrb1/M11_d
+ N_C[10]_XADDER/Xa011/Xrb1/M11_g N_VDD_XADDER/Xa011/Xrb1/M11_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXBOOTH/Xsel26/M14 N_PP2[6]_XBOOTH/Xsel26/M14_d
+ N_XBOOTH/XSEL26/N004_XBOOTH/Xsel26/M14_g N_VDD_XBOOTH/Xsel26/M14_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel16/M14 N_PP1[6]_XBOOTH/Xsel16/M14_d
+ N_XBOOTH/XSEL16/N004_XBOOTH/Xsel16/M14_g N_VDD_XBOOTH/Xsel16/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXBOOTH/Xsel06/M14 N_PP0[6]_XBOOTH/Xsel06/M14_d
+ N_XBOOTH/XSEL06/N004_XBOOTH/Xsel06/M14_g N_VDD_XBOOTH/Xsel06/M14_s
+ N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/X_LV3_FA10/M28 N_XCSA/LV3_C[13]_XCSA/X_LV3_FA10/M28_d
+ N_XCSA/X_LV3_FA10/_COUT_XCSA/X_LV3_FA10/M28_g N_VDD_XCSA/X_LV3_FA10/M28_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXADDER/Xa710/M4 N_OUT1[10]_XADDER/Xa710/M4_d
+ N_XADDER/XA710/N002_XADDER/Xa710/M4_g N_VDD_XADDER/Xa710/M4_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa712/M5 N_XADDER/XA712/N002_XADDER/Xa712/M5_d
+ N_XADDER/P12_XADDER/Xa712/M5_g N_XADDER/XA712/N001_XADDER/Xa712/M5_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=4.444e-13 AS=6.16e-14
+ PD=2.46e-06 PS=2.8e-07
mX02/xd212/M4 N_X02/XD212/N1_X02/xd212/M4_d N_CLK_X02/xd212/M4_g
+ N_VDD_X02/xd212/M4_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA9/M28 N_XCSA/LV3_C[12]_XCSA/X_LV3_FA9/M28_d
+ N_XCSA/X_LV3_FA9/_COUT_XCSA/X_LV3_FA9/M28_g N_VDD_XCSA/X_LV3_FA9/M28_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXCSA/Xdffa10/M4 N_XCSA/XDFFA10/N1_XCSA/Xdffa10/M4_d N_CLK_XCSA/Xdffa10/M4_g
+ N_VDD_XCSA/Xdffa10/M4_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa23/M4 N_XCSA/XDFFA23/N1_XCSA/Xdffa23/M4_d N_CLK_XCSA/Xdffa23/M4_g
+ N_VDD_XCSA/Xdffa23/M4_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA10/M27 N_XCSA/LV3_S[12]_XCSA/X_LV3_FA10/M27_d
+ N_XCSA/X_LV3_FA10/_SUM_XCSA/X_LV3_FA10/M27_g N_VDD_XCSA/X_LV3_FA10/M27_s
+ N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mX02/xd212/M7 N_X02/XD212/N3_X02/xd212/M7_d N_X02/XD212/N1_X02/xd212/M7_g
+ N_VDD_X02/xd212/M7_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/X_LV3_FA9/M27 N_XCSA/LV3_S[11]_XCSA/X_LV3_FA9/M27_d
+ N_XCSA/X_LV3_FA9/_SUM_XCSA/X_LV3_FA9/M27_g N_VDD_XCSA/X_LV3_FA9/M27_s
+ N_VDD_XACCXOR/X_xor2/M4_b P_18_G2 L=1.8e-07 W=5.5e-07 AD=2.695e-13 AS=2.695e-13
+ PD=1.53e-06 PS=1.53e-06
mXCSA/Xdffa10/M7 N_XCSA/XDFFA10/N3_XCSA/Xdffa10/M7_d
+ N_XCSA/XDFFA10/N1_XCSA/Xdffa10/M7_g N_VDD_XCSA/Xdffa10/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa23/M7 N_XCSA/XDFFA23/N3_XCSA/Xdffa23/M7_d
+ N_XCSA/XDFFA23/N1_XCSA/Xdffa23/M7_g N_VDD_XCSA/Xdffa23/M7_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa011/Xrb1/Xand1/M15 N_VDD_XADDER/Xa011/Xrb1/Xand1/M15_d
+ N_XADDER/XA011/XRB1/N003_XADDER/Xa011/Xrb1/Xand1/M15_g
+ N_XADDER/G10_XADDER/Xa011/Xrb1/Xand1/M15_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/X_inv2/mp N_XCSA/PP2_INVS_XCSA/X_inv2/mp_d N_PP2[6]_XCSA/X_inv2/mp_g
+ N_VDD_XCSA/X_inv2/mp_s N_VDD_XBOOTH/Xdffa4/M1_b P_18_G2 L=1.8e-07 W=5.5e-07
+ AD=2.695e-13 AS=2.695e-13 PD=1.53e-06 PS=1.53e-06
mXCSA/X_inv1/mp N_XCSA/PP1_INVS_XCSA/X_inv1/mp_d N_PP1[6]_XCSA/X_inv1/mp_g
+ N_VDD_XCSA/X_inv1/mp_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=5.5e-07
+ AD=2.695e-13 AS=2.695e-13 PD=1.53e-06 PS=1.53e-06
mXCSA/X_inv0/mp N_XCSA/PP0_INVS_XCSA/X_inv0/mp_d N_PP0[6]_XCSA/X_inv0/mp_g
+ N_VDD_XCSA/X_inv0/mp_s N_VDD_XBOOTH/Xdffa2/M1_b P_18_G2 L=1.8e-07 W=5.5e-07
+ AD=2.695e-13 AS=2.695e-13 PD=1.53e-06 PS=1.53e-06
mXADDER/Xa111/Xyb1/M11 N_XADDER/XA111/XYB1/N003_XADDER/Xa111/Xyb1/M11_d
+ N_XADDER/P10_XADDER/Xa111/Xyb1/M11_g N_VDD_XADDER/Xa111/Xyb1/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mXADDER/Xa710/M5 N_XADDER/XA710/N002_XADDER/Xa710/M5_d
+ N_XADDER/P10_XADDER/Xa710/M5_g N_XADDER/XA710/N001_XADDER/Xa710/M5_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=4.444e-13 AS=6.16e-14
+ PD=2.46e-06 PS=2.8e-07
mXADDER/Xa712/M4 N_OUT1[12]_XADDER/Xa712/M4_d
+ N_XADDER/XA712/N002_XADDER/Xa712/M4_g N_VDD_XADDER/Xa712/M4_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa111/Xyb1/M12 N_XADDER/XA111/XYB1/N003_XADDER/Xa111/Xyb1/M12_d
+ N_XADDER/P11_XADDER/Xa111/Xyb1/M12_g N_VDD_XADDER/Xa111/Xyb1/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd212/M10 N_OUT[11]_X02/xd212/M10_d N_X02/XD212/N3_X02/xd212/M10_g
+ N_VDD_X02/xd212/M10_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa710/M6 N_XADDER/XA710/N001_XADDER/Xa710/M6_d
+ N_XADDER/GX5[1]_XADDER/Xa710/M6_g N_VDD_XADDER/Xa710/M6_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa10/M10 N_C[11]_XCSA/Xdffa10/M10_d
+ N_XCSA/XDFFA10/N3_XCSA/Xdffa10/M10_g N_VDD_XCSA/Xdffa10/M10_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa23/M10 N_S[11]_XCSA/Xdffa23/M10_d
+ N_XCSA/XDFFA23/N3_XCSA/Xdffa23/M10_g N_VDD_XCSA/Xdffa23/M10_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa012/Xrb2/M4 N_XADDER/P11_XADDER/Xa012/Xrb2/M4_d
+ N_XADDER/XA012/XRB2/N002_XADDER/Xa012/Xrb2/M4_g N_VDD_XADDER/Xa012/Xrb2/M4_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa111/Xyb2/M12 N_XADDER/XA111/XYB2/N003_XADDER/Xa111/Xyb2/M12_d
+ N_XADDER/P11_XADDER/Xa111/Xyb2/M12_g N_VDD_XADDER/Xa111/Xyb2/M12_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mX02/xd213/M1 N_X02/XD213/P001_X02/xd213/M1_d N_OUT1[12]_X02/xd213/M1_g
+ N_VDD_X02/xd213/M1_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14
+ AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXADDER/Xa013/M6 N_XADDER/XA013/N001_XADDER/Xa013/M6_d N_C[12]_XADDER/Xa013/M6_g
+ N_VDD_XADDER/Xa013/M6_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=6.16e-14 AS=2.156e-13 PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa11/M1 N_XCSA/XDFFA11/P001_XCSA/Xdffa11/M1_d
+ N_XCSA/LV3_C[12]_XCSA/Xdffa11/M1_g N_VDD_XCSA/Xdffa11/M1_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXCSA/Xdffa24/M1 N_XCSA/XDFFA24/P001_XCSA/Xdffa24/M1_d
+ N_XCSA/LV3_S[12]_XCSA/Xdffa24/M1_g N_VDD_XCSA/Xdffa24/M1_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXADDER/Xa111/Xyb2/M11 N_XADDER/XA111/XYB2/N003_XADDER/Xa111/Xyb2/M11_d
+ N_XADDER/G10_XADDER/Xa111/Xyb2/M11_g N_VDD_XADDER/Xa111/Xyb2/M11_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.86e-13 AS=1.188e-13
+ PD=1.74e-06 PS=5.4e-07
mX02/xd213/M2 N_X02/XD213/N0_X02/xd213/M2_d N_CLK_X02/xd213/M2_g
+ N_X02/XD213/P001_X02/xd213/M2_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa012/Xrb2/M5 N_XADDER/XA012/XRB2/N001_XADDER/Xa012/Xrb2/M5_d
+ N_C[11]_XADDER/Xa012/Xrb2/M5_g N_VDD_XADDER/Xa012/Xrb2/M5_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.904e-13
+ PD=2.8e-07 PS=1.76e-06
mXADDER/Xa013/M5 N_XADDER/XA013/N002_XADDER/Xa013/M5_d N_S[12]_XADDER/Xa013/M5_g
+ N_XADDER/XA013/N001_XADDER/Xa013/M5_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=4.444e-13 AS=6.16e-14 PD=2.46e-06 PS=2.8e-07
mXCSA/Xdffa11/M2 N_XCSA/XDFFA11/N0_XCSA/Xdffa11/M2_d N_CLK_XCSA/Xdffa11/M2_g
+ N_XCSA/XDFFA11/P001_XCSA/Xdffa11/M2_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXCSA/Xdffa24/M2 N_XCSA/XDFFA24/N0_XCSA/Xdffa24/M2_d N_CLK_XCSA/Xdffa24/M2_g
+ N_XCSA/XDFFA24/P001_XCSA/Xdffa24/M2_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07
+ W=4.4e-07 AD=2.156e-13 AS=6.16e-14 PD=1.42e-06 PS=2.8e-07
mXADDER/Xa711/M4 N_OUT1[11]_XADDER/Xa711/M4_d
+ N_XADDER/XA711/N002_XADDER/Xa711/M4_g N_VDD_XADDER/Xa711/M4_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa012/Xrb2/M6 N_XADDER/XA012/XRB2/N002_XADDER/Xa012/Xrb2/M6_d
+ N_S[11]_XADDER/Xa012/Xrb2/M6_g N_XADDER/XA012/XRB2/N001_XADDER/Xa012/Xrb2/M6_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=6.16e-14
+ PD=1.42e-06 PS=2.8e-07
mX02/xd213/M4 N_X02/XD213/N1_X02/xd213/M4_d N_CLK_X02/xd213/M4_g
+ N_VDD_X02/xd213/M4_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXADDER/Xa111/Xyb2/Xand1/M15 N_VDD_XADDER/Xa111/Xyb2/Xand1/M15_d
+ N_XADDER/XA111/XYB2/N003_XADDER/Xa111/Xyb2/Xand1/M15_g
+ N_XADDER/XA111/T1_XADDER/Xa111/Xyb2/Xand1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa11/M4 N_XCSA/XDFFA11/N1_XCSA/Xdffa11/M4_d N_CLK_XCSA/Xdffa11/M4_g
+ N_VDD_XCSA/Xdffa11/M4_s N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa24/M4 N_XCSA/XDFFA24/N1_XCSA/Xdffa24/M4_d N_CLK_XCSA/Xdffa24/M4_g
+ N_VDD_XCSA/Xdffa24/M4_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mX02/xd213/M7 N_X02/XD213/N3_X02/xd213/M7_d N_X02/XD213/N1_X02/xd213/M7_g
+ N_VDD_X02/xd213/M7_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13
+ AS=1.188e-13 PD=1.42e-06 PS=5.4e-07
mXADDER/Xa013/M4 N_XADDER/P12_XADDER/Xa013/M4_d
+ N_XADDER/XA013/N002_XADDER/Xa013/M4_g N_VDD_XADDER/Xa013/M4_s
+ N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa012/Xrb1/M12 N_XADDER/XA012/XRB1/N003_XADDER/Xa012/Xrb1/M12_d
+ N_S[11]_XADDER/Xa012/Xrb1/M12_g N_VDD_XADDER/Xa012/Xrb1/M12_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa711/M5 N_XADDER/XA711/N002_XADDER/Xa711/M5_d
+ N_XADDER/P11_XADDER/Xa711/M5_g N_XADDER/XA711/N001_XADDER/Xa711/M5_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=4.444e-13 AS=6.16e-14
+ PD=2.46e-06 PS=2.8e-07
mXCSA/Xdffa11/M7 N_XCSA/XDFFA11/N3_XCSA/Xdffa11/M7_d
+ N_XCSA/XDFFA11/N1_XCSA/Xdffa11/M7_g N_VDD_XCSA/Xdffa11/M7_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXCSA/Xdffa24/M7 N_XCSA/XDFFA24/N3_XCSA/Xdffa24/M7_d
+ N_XCSA/XDFFA24/N1_XCSA/Xdffa24/M7_g N_VDD_XCSA/Xdffa24/M7_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa711/M6 N_XADDER/XA711/N001_XADDER/Xa711/M6_d
+ N_XADDER/GX6[4]_XADDER/Xa711/M6_g N_VDD_XADDER/Xa711/M6_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=6.16e-14 AS=2.156e-13
+ PD=2.8e-07 PS=1.42e-06
mXADDER/Xa012/Xrb1/M11 N_XADDER/XA012/XRB1/N003_XADDER/Xa012/Xrb1/M11_d
+ N_C[11]_XADDER/Xa012/Xrb1/M11_g N_VDD_XADDER/Xa012/Xrb1/M11_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.188e-13
+ PD=1.42e-06 PS=5.4e-07
mXADDER/Xa111/Xyb3/M36 N_XADDER/XA111/XYB3/N008_XADDER/Xa111/Xyb3/M36_d
+ N_XADDER/XA111/T1_XADDER/Xa111/Xyb3/M36_g
+ N_XADDER/XA111/XYB3/N007_XADDER/Xa111/Xyb3/M36_s N_VDD_XADDER/Xa000/Xao1/M12_b
+ P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=1.21e-13 PD=1.42e-06 PS=5.5e-07
mX02/xd213/M10 N_OUT[12]_X02/xd213/M10_d N_X02/XD213/N3_X02/xd213/M10_g
+ N_VDD_X02/xd213/M10_s N_VDD_XADDER/Xa72/M4_b P_18_G2 L=1.8e-07 W=4.4e-07
+ AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa111/Xyb3/M35 N_XADDER/XA111/XYB3/N007_XADDER/Xa111/Xyb3/M35_d
+ N_XADDER/G11_XADDER/Xa111/Xyb3/M35_g N_VDD_XADDER/Xa111/Xyb3/M35_s
+ N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=1.21e-13 AS=1.298e-13
+ PD=5.5e-07 PS=5.9e-07
mXCSA/Xdffa11/M10 N_C[12]_XCSA/Xdffa11/M10_d
+ N_XCSA/XDFFA11/N3_XCSA/Xdffa11/M10_g N_VDD_XCSA/Xdffa11/M10_s
+ N_VDD_XACCXOR/X_xor1/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXCSA/Xdffa24/M10 N_S[12]_XCSA/Xdffa24/M10_d
+ N_XCSA/XDFFA24/N3_XCSA/Xdffa24/M10_g N_VDD_XCSA/Xdffa24/M10_s
+ N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2 L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13
+ PD=1.42e-06 PS=1.42e-06
mXADDER/Xa012/Xrb1/Xand1/M15 N_VDD_XADDER/Xa012/Xrb1/Xand1/M15_d
+ N_XADDER/XA012/XRB1/N003_XADDER/Xa012/Xrb1/Xand1/M15_g
+ N_XADDER/G11_XADDER/Xa012/Xrb1/Xand1/M15_s N_VDD_XADDER/Xa01/Xrb2/M4_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=2.156e-13 AS=2.156e-13 PD=1.42e-06 PS=1.42e-06
mXADDER/Xa111/Xyb3/Xor1/M15 N_VDD_XADDER/Xa111/Xyb3/Xor1/M15_d
+ N_XADDER/XA111/XYB3/N008_XADDER/Xa111/Xyb3/Xor1/M15_g
+ N_XADDER/GG11_XADDER/Xa111/Xyb3/Xor1/M15_s N_VDD_XADDER/Xa000/Xao1/M12_b P_18_G2
+ L=1.8e-07 W=4.4e-07 AD=1.298e-13 AS=3.916e-13 PD=5.9e-07 PS=2.22e-06
*
.include "MAC6_LPE.sp.MAC6.pxi"
*
.ends
*
*
